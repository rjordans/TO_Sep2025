magic
tech ihp-sg13g2
magscale 1 2
timestamp 1756455342
<< nwell >>
rect -1596 1288 183 2631
rect -1596 1028 -939 1288
rect -1596 813 -1136 1028
<< hvnmos >>
rect -1320 528 -1260 618
rect -1033 528 -973 618
rect -1320 362 -1260 452
rect -688 686 -288 1086
rect -194 686 206 1086
rect -688 86 -288 486
rect -194 86 206 486
<< hvpmos >>
rect -1320 1961 -1260 2361
rect -1320 1483 -1260 1883
rect -987 2196 -587 2296
rect -511 2196 -111 2296
rect -987 2008 -587 2108
rect -511 2008 -111 2108
rect -987 1820 -587 1920
rect -511 1820 -111 1920
rect -987 1632 -587 1732
rect -511 1632 -111 1732
rect -1320 1005 -1260 1405
rect -1129 1221 -1069 1301
<< hvndiff >>
rect -688 1141 -288 1155
rect -688 1108 -674 1141
rect -307 1108 -288 1141
rect -688 1086 -288 1108
rect -194 1149 206 1163
rect -194 1116 -180 1149
rect 187 1116 206 1149
rect -194 1086 206 1116
rect -1320 672 -1260 689
rect -1320 640 -1306 672
rect -1274 640 -1260 672
rect -1320 618 -1260 640
rect -1033 672 -973 689
rect -1033 640 -1019 672
rect -987 640 -973 672
rect -1033 618 -973 640
rect -1320 506 -1260 528
rect -1320 474 -1306 506
rect -1274 474 -1260 506
rect -1320 452 -1260 474
rect -1033 506 -973 528
rect -1033 474 -1019 506
rect -987 474 -973 506
rect -1033 460 -973 474
rect -1320 340 -1260 362
rect -1320 307 -1306 340
rect -1274 307 -1260 340
rect -1320 293 -1260 307
rect -688 656 -288 686
rect -688 623 -669 656
rect -302 623 -288 656
rect -688 605 -288 623
rect -194 652 206 686
rect -194 619 -180 652
rect 187 619 206 652
rect -688 549 -288 563
rect -688 516 -674 549
rect -307 516 -288 549
rect -688 486 -288 516
rect -194 549 206 619
rect -194 516 -180 549
rect 187 516 206 549
rect -194 486 206 516
rect -688 52 -288 86
rect -688 19 -669 52
rect -302 19 -288 52
rect -688 5 -288 19
rect -194 52 206 86
rect -194 19 -180 52
rect 187 19 206 52
rect -194 5 206 19
<< hvpdiff >>
rect -1320 2423 -1260 2441
rect -1320 2391 -1306 2423
rect -1274 2391 -1260 2423
rect -1320 2361 -1260 2391
rect -1320 1939 -1260 1961
rect -1320 1907 -1306 1939
rect -1274 1907 -1260 1939
rect -1320 1883 -1260 1907
rect -1320 1461 -1260 1483
rect -1320 1429 -1306 1461
rect -1274 1429 -1260 1461
rect -1320 1405 -1260 1429
rect -1055 2282 -987 2296
rect -1055 2210 -1041 2282
rect -1009 2210 -987 2282
rect -1055 2196 -987 2210
rect -587 2282 -511 2296
rect -587 2210 -565 2282
rect -533 2210 -511 2282
rect -587 2196 -511 2210
rect -111 2282 -43 2296
rect -111 2210 -89 2282
rect -57 2210 -43 2282
rect -111 2196 -43 2210
rect -1055 2094 -987 2108
rect -1055 2022 -1041 2094
rect -1009 2022 -987 2094
rect -1055 2008 -987 2022
rect -587 2094 -511 2108
rect -587 2022 -565 2094
rect -533 2022 -511 2094
rect -587 2008 -511 2022
rect -111 2094 -43 2108
rect -111 2022 -89 2094
rect -57 2022 -43 2094
rect -111 2008 -43 2022
rect -1055 1906 -987 1920
rect -1055 1834 -1041 1906
rect -1009 1834 -987 1906
rect -1055 1820 -987 1834
rect -587 1906 -511 1920
rect -587 1834 -565 1906
rect -533 1834 -511 1906
rect -587 1820 -511 1834
rect -111 1906 -43 1920
rect -111 1834 -89 1906
rect -57 1834 -43 1906
rect -111 1820 -43 1834
rect -1055 1718 -987 1732
rect -1055 1646 -1041 1718
rect -1009 1646 -987 1718
rect -1055 1632 -987 1646
rect -587 1718 -511 1732
rect -587 1646 -565 1718
rect -533 1646 -511 1718
rect -587 1632 -511 1646
rect -111 1718 -43 1732
rect -111 1646 -89 1718
rect -57 1646 -43 1718
rect -111 1632 -43 1646
rect -1129 1355 -1069 1369
rect -1129 1323 -1115 1355
rect -1083 1323 -1069 1355
rect -1129 1301 -1069 1323
rect -1129 1199 -1069 1221
rect -1129 1167 -1115 1199
rect -1083 1167 -1069 1199
rect -1129 1153 -1069 1167
rect -1320 983 -1260 1005
rect -1320 951 -1306 983
rect -1274 951 -1260 983
rect -1320 937 -1260 951
<< hvndiffc >>
rect -674 1108 -307 1141
rect -180 1116 187 1149
rect -1306 640 -1274 672
rect -1019 640 -987 672
rect -1306 474 -1274 506
rect -1019 474 -987 506
rect -1306 307 -1274 340
rect -669 623 -302 656
rect -180 619 187 652
rect -674 516 -307 549
rect -180 516 187 549
rect -669 19 -302 52
rect -180 19 187 52
<< hvpdiffc >>
rect -1306 2391 -1274 2423
rect -1306 1907 -1274 1939
rect -1306 1429 -1274 1461
rect -1041 2210 -1009 2282
rect -565 2210 -533 2282
rect -89 2210 -57 2282
rect -1041 2022 -1009 2094
rect -565 2022 -533 2094
rect -89 2022 -57 2094
rect -1041 1834 -1009 1906
rect -565 1834 -533 1906
rect -89 1834 -57 1906
rect -1041 1646 -1009 1718
rect -565 1646 -533 1718
rect -89 1646 -57 1718
rect -1115 1323 -1083 1355
rect -1115 1167 -1083 1199
rect -1306 951 -1274 983
<< psubdiff >>
rect 320 2365 1820 2379
rect 320 29 334 2365
rect 366 2319 1774 2333
rect 366 75 380 2319
rect 1760 75 1774 2319
rect 366 61 1774 75
rect 1806 29 1820 2365
rect 320 15 1820 29
<< hvpsubdiff >>
rect -870 868 -810 882
rect -1472 639 -1412 653
rect -1472 113 -1458 639
rect -1426 159 -1412 639
rect -870 159 -856 868
rect -1426 145 -856 159
rect -902 113 -856 145
rect -824 113 -810 868
rect -1472 99 -810 113
<< hvnsubdiff >>
rect -1472 2493 -1260 2507
rect -1472 951 -1458 2493
rect -1274 2461 -1260 2493
rect -1426 2447 -1260 2461
rect -1426 951 -1412 2447
rect -1320 2441 -1260 2447
rect -1157 2493 59 2507
rect -1157 1426 -1143 2493
rect -1111 2447 13 2461
rect -1111 1472 -1097 2447
rect -1 1472 13 2447
rect -1111 1458 13 1472
rect 45 1426 59 2493
rect -1157 1412 59 1426
rect -1472 937 -1412 951
<< psubdiffcont >>
rect 334 2333 1806 2365
rect 334 61 366 2333
rect 1774 61 1806 2333
rect 334 29 1806 61
<< hvpsubdiffcont >>
rect -1458 145 -1426 639
rect -1458 113 -902 145
rect -856 113 -824 868
<< hvnsubdiffcont >>
rect -1458 2461 -1274 2493
rect -1458 951 -1426 2461
rect -1143 2461 45 2493
rect -1143 1458 -1111 2461
rect 13 1458 45 2461
rect -1143 1426 45 1458
<< poly >>
rect -1394 2339 -1320 2361
rect -1394 1981 -1380 2339
rect -1348 1981 -1320 2339
rect -1394 1961 -1320 1981
rect -1260 1961 -1212 2361
rect -1394 1861 -1320 1883
rect -1394 1503 -1380 1861
rect -1348 1503 -1320 1861
rect -1394 1483 -1320 1503
rect -1260 1483 -1212 1883
rect -987 2356 -587 2374
rect -987 2324 -973 2356
rect -609 2324 -587 2356
rect -987 2296 -587 2324
rect -511 2356 -111 2374
rect -511 2324 -489 2356
rect -125 2324 -111 2356
rect -511 2296 -111 2324
rect -987 2168 -587 2196
rect -987 2136 -973 2168
rect -609 2136 -587 2168
rect -987 2108 -587 2136
rect -511 2168 -111 2196
rect -511 2136 -489 2168
rect -125 2136 -111 2168
rect -511 2108 -111 2136
rect -987 1980 -587 2008
rect -987 1948 -973 1980
rect -609 1948 -587 1980
rect -987 1920 -587 1948
rect -511 1980 -111 2008
rect -511 1948 -489 1980
rect -125 1948 -111 1980
rect -511 1920 -111 1948
rect -987 1792 -587 1820
rect -987 1760 -973 1792
rect -609 1760 -587 1792
rect -987 1732 -587 1760
rect -511 1792 -111 1820
rect -511 1760 -489 1792
rect -125 1760 -111 1792
rect -511 1732 -111 1760
rect -987 1604 -587 1632
rect -987 1572 -973 1604
rect -609 1572 -587 1604
rect -987 1558 -587 1572
rect -511 1604 -111 1632
rect -511 1572 -489 1604
rect -125 1572 -111 1604
rect -511 1558 -111 1572
rect -1394 1383 -1320 1405
rect -1394 1025 -1380 1383
rect -1348 1025 -1320 1383
rect -1394 1005 -1320 1025
rect -1260 1005 -1212 1405
rect -1176 1221 -1129 1301
rect -1069 1278 -985 1301
rect -1069 1246 -1034 1278
rect -1002 1246 -985 1278
rect -1069 1221 -985 1246
rect -770 1072 -688 1086
rect -1395 604 -1320 618
rect -1395 542 -1380 604
rect -1348 542 -1320 604
rect -1395 528 -1320 542
rect -1260 528 -1214 618
rect -1079 528 -1033 618
rect -973 604 -898 618
rect -973 542 -945 604
rect -912 542 -898 604
rect -973 528 -898 542
rect -1366 362 -1320 452
rect -1260 438 -1185 452
rect -1260 376 -1232 438
rect -1200 376 -1185 438
rect -1260 362 -1185 376
rect -770 700 -748 1072
rect -716 700 -688 1072
rect -770 686 -688 700
rect -288 1072 -194 1086
rect -288 700 -260 1072
rect -222 700 -194 1072
rect -288 686 -194 700
rect 206 1072 280 1086
rect 206 700 234 1072
rect 266 700 280 1072
rect 206 686 280 700
rect -770 472 -688 486
rect -770 100 -748 472
rect -716 100 -688 472
rect -770 86 -688 100
rect -288 472 -194 486
rect -288 100 -260 472
rect -222 100 -194 472
rect -288 86 -194 100
rect 206 472 280 486
rect 206 100 234 472
rect 266 100 280 472
rect 206 86 280 100
rect 460 2269 560 2283
rect 460 2237 474 2269
rect 546 2237 560 2269
rect 460 2197 560 2237
rect 460 157 560 197
rect 460 125 474 157
rect 546 125 560 157
rect 460 111 560 125
rect 620 2269 720 2283
rect 620 2237 634 2269
rect 706 2237 720 2269
rect 620 2197 720 2237
rect 620 157 720 197
rect 620 125 634 157
rect 706 125 720 157
rect 620 110 720 125
rect 780 2269 880 2283
rect 780 2237 794 2269
rect 866 2237 880 2269
rect 780 2197 880 2237
rect 780 157 880 197
rect 780 125 794 157
rect 866 125 880 157
rect 780 110 880 125
rect 940 2269 1040 2283
rect 940 2237 954 2269
rect 1026 2237 1040 2269
rect 940 2197 1040 2237
rect 940 157 1040 197
rect 940 125 954 157
rect 1026 125 1040 157
rect 940 110 1040 125
rect 1100 2269 1200 2283
rect 1100 2237 1114 2269
rect 1186 2237 1200 2269
rect 1100 2197 1200 2237
rect 1100 157 1200 197
rect 1100 125 1114 157
rect 1186 125 1200 157
rect 1100 110 1200 125
rect 1260 2269 1360 2283
rect 1260 2237 1274 2269
rect 1346 2237 1360 2269
rect 1260 2197 1360 2237
rect 1260 157 1360 197
rect 1260 125 1274 157
rect 1346 125 1360 157
rect 1260 110 1360 125
rect 1420 2269 1520 2283
rect 1420 2237 1434 2269
rect 1506 2237 1520 2269
rect 1420 2197 1520 2237
rect 1420 157 1520 197
rect 1420 125 1434 157
rect 1506 125 1520 157
rect 1420 110 1520 125
rect 1580 2269 1680 2283
rect 1580 2237 1594 2269
rect 1666 2237 1680 2269
rect 1580 2197 1680 2237
rect 1580 157 1680 197
rect 1580 125 1594 157
rect 1666 125 1680 157
rect 1580 110 1680 125
<< polycont >>
rect -1380 1981 -1348 2339
rect -1380 1503 -1348 1861
rect -973 2324 -609 2356
rect -489 2324 -125 2356
rect -973 2136 -609 2168
rect -489 2136 -125 2168
rect -973 1948 -609 1980
rect -489 1948 -125 1980
rect -973 1760 -609 1792
rect -489 1760 -125 1792
rect -973 1572 -609 1604
rect -489 1572 -125 1604
rect -1380 1025 -1348 1383
rect -1034 1246 -1002 1278
rect -1380 542 -1348 604
rect -945 542 -912 604
rect -1232 376 -1200 438
rect -748 700 -716 1072
rect -260 700 -222 1072
rect 234 700 266 1072
rect -748 100 -716 472
rect -260 100 -222 472
rect 234 100 266 472
rect 474 2237 546 2269
rect 474 125 546 157
rect 634 2237 706 2269
rect 634 125 706 157
rect 794 2237 866 2269
rect 794 125 866 157
rect 954 2237 1026 2269
rect 954 125 1026 157
rect 1114 2237 1186 2269
rect 1114 125 1186 157
rect 1274 2237 1346 2269
rect 1274 125 1346 157
rect 1434 2237 1506 2269
rect 1434 125 1506 157
rect 1594 2237 1666 2269
rect 1594 125 1666 157
<< ppolyres >>
rect 460 197 560 2197
rect 620 197 720 2197
rect 780 197 880 2197
rect 940 197 1040 2197
rect 1100 197 1200 2197
rect 1260 197 1360 2197
rect 1420 197 1520 2197
rect 1580 197 1680 2197
<< metal1 >>
rect -1468 2493 55 2503
rect -1468 951 -1458 2493
rect -1274 2461 -1143 2493
rect -1426 2451 -1143 2461
rect -1426 951 -1416 2451
rect -1306 2423 -1274 2451
rect -1306 2381 -1274 2391
rect -1153 2365 -1143 2451
rect -1111 2451 13 2461
rect -1380 2339 -1348 2349
rect -1380 1939 -1348 1981
rect -1380 1907 -1306 1939
rect -1274 1907 -1264 1939
rect -1380 1861 -1348 1871
rect -1380 1461 -1348 1503
rect -1380 1429 -1306 1461
rect -1274 1429 -1264 1461
rect -1153 1425 -1152 2365
rect -1111 1468 -1103 2451
rect -973 2356 -609 2367
rect -1057 2282 -1009 2296
rect -1057 2206 -1053 2282
rect -1013 2206 -1009 2210
rect -1057 2197 -1009 2206
rect -973 2168 -965 2324
rect -620 2168 -609 2324
rect -973 2104 -965 2136
rect -1041 2094 -965 2104
rect -1009 2022 -965 2094
rect -1041 2012 -965 2022
rect -973 1987 -965 2012
rect -620 1987 -609 2136
rect -973 1980 -609 1987
rect -1060 1908 -1009 1920
rect -1060 1836 -1050 1908
rect -1010 1906 -1009 1908
rect -1060 1834 -1041 1836
rect -1060 1824 -1009 1834
rect -973 1792 -609 1948
rect -1060 1721 -1009 1732
rect -1060 1645 -1055 1721
rect -1015 1718 -1009 1721
rect -1015 1645 -1009 1646
rect -1060 1636 -1009 1645
rect -973 1604 -609 1760
rect -973 1561 -609 1572
rect -565 2282 -533 2451
rect -565 2094 -533 2210
rect -565 1906 -533 2022
rect -565 1718 -533 1834
rect -565 1468 -533 1646
rect -489 2356 -125 2366
rect -489 2168 -482 2324
rect -155 2182 -125 2324
rect -89 2284 -46 2296
rect -89 2282 -87 2284
rect -89 2208 -87 2210
rect -47 2208 -46 2284
rect -89 2197 -46 2208
rect -320 2168 -125 2182
rect -489 1986 -482 2136
rect -320 1986 -125 2136
rect -89 2094 -47 2105
rect -48 2022 -47 2094
rect -89 2012 -47 2022
rect -489 1980 -125 1986
rect -489 1917 -125 1948
rect -489 1906 -47 1917
rect -489 1834 -89 1906
rect -57 1834 -47 1906
rect -489 1824 -47 1834
rect -489 1792 -125 1824
rect -489 1604 -475 1760
rect -143 1604 -125 1760
rect -89 1718 -47 1729
rect -48 1646 -47 1718
rect -89 1636 -47 1646
rect -489 1561 -125 1572
rect 5 1468 13 2451
rect -1111 1458 13 1468
rect 45 1426 55 2493
rect -1112 1425 55 1426
rect -1153 1416 55 1425
rect 324 2373 1816 2375
rect 324 2365 413 2373
rect 1798 2365 1816 2373
rect 324 2364 334 2365
rect -1468 941 -1416 951
rect -1380 1383 -1348 1393
rect -1126 1355 -1073 1416
rect -1126 1323 -1115 1355
rect -1083 1323 -1073 1355
rect -522 1346 -281 1359
rect -522 1344 -509 1346
rect -1126 1313 -1073 1323
rect -1036 1322 -509 1344
rect -1037 1308 -509 1322
rect -1037 1278 -1001 1308
rect -522 1306 -509 1308
rect -296 1344 -281 1346
rect -100 1346 -42 1347
rect -100 1344 -91 1346
rect -296 1308 -91 1344
rect -296 1306 -281 1308
rect -522 1296 -281 1306
rect -100 1306 -91 1308
rect -51 1306 -42 1346
rect -100 1305 -42 1306
rect -1037 1246 -1034 1278
rect -1002 1246 -1001 1278
rect 324 1252 331 2364
rect -1380 885 -1348 1025
rect -1130 1199 -1078 1209
rect -1130 1167 -1115 1199
rect -1083 1167 -1078 1199
rect -1130 1091 -1078 1167
rect -1439 873 -1348 885
rect -1439 721 -1430 873
rect -1359 721 -1348 873
rect -1439 708 -1348 721
rect -1468 639 -1416 649
rect -1468 113 -1458 639
rect -1426 155 -1416 639
rect -1380 604 -1348 708
rect -1306 983 -1274 994
rect -1306 884 -1274 951
rect -1130 991 -1079 1091
rect -1037 1078 -1001 1246
rect -866 1200 331 1252
rect -1037 1042 -909 1078
rect -1130 974 -997 991
rect -1306 875 -1241 884
rect -1306 768 -1293 875
rect -1253 768 -1241 875
rect -1306 756 -1241 768
rect -1306 705 -1274 756
rect -1306 672 -1255 705
rect -1274 640 -1255 672
rect -1306 630 -1255 640
rect -1130 661 -1105 974
rect -1023 684 -997 974
rect -1023 672 -987 684
rect -1023 661 -1019 672
rect -1130 640 -1019 661
rect -1130 630 -987 640
rect -945 604 -909 1042
rect -866 868 -814 1200
rect -191 1157 197 1158
rect -191 1149 -179 1157
rect -685 1108 -674 1141
rect -307 1108 -297 1141
rect -191 1116 -180 1149
rect 188 1117 197 1157
rect 187 1116 197 1117
rect -685 1072 -297 1108
rect -955 542 -945 604
rect -912 542 -902 604
rect -1380 530 -1348 542
rect -1033 506 -981 507
rect -866 506 -856 868
rect -1320 474 -1306 506
rect -1274 474 -1019 506
rect -987 474 -856 506
rect -1033 460 -945 474
rect -1301 429 -1232 438
rect -1301 384 -1292 429
rect -1301 376 -1232 384
rect -1200 376 -1189 438
rect -1316 329 -1306 340
rect -1274 329 -1264 340
rect -1316 257 -1310 329
rect -1270 257 -1264 329
rect -1316 248 -1264 257
rect -866 155 -856 474
rect -1426 145 -856 155
rect -902 113 -856 145
rect -824 656 -814 868
rect -770 700 -748 1072
rect -716 1046 -260 1072
rect -333 713 -260 1046
rect -716 700 -260 713
rect -222 700 234 1072
rect 266 700 280 1072
rect 324 692 331 1200
rect 371 2325 413 2333
rect 371 2323 1774 2325
rect 371 692 376 2323
rect 463 2269 716 2279
rect 463 2237 474 2269
rect 546 2237 634 2269
rect 706 2237 716 2269
rect 463 2227 716 2237
rect 783 2269 1036 2279
rect 783 2237 794 2269
rect 866 2237 954 2269
rect 1026 2237 1036 2269
rect 783 2227 1036 2237
rect 1103 2269 1356 2279
rect 1103 2237 1114 2269
rect 1186 2237 1274 2269
rect 1346 2237 1356 2269
rect 1103 2227 1356 2237
rect 1423 2269 1676 2279
rect 1423 2237 1434 2269
rect 1506 2237 1594 2269
rect 1666 2237 1676 2269
rect 1423 2227 1676 2237
rect 1764 2268 1774 2323
rect 1806 2268 1816 2365
rect -824 623 -669 656
rect -302 623 -292 656
rect -192 652 198 656
rect -824 508 -721 623
rect -192 619 -180 652
rect 187 619 198 652
rect -192 549 31 619
rect 184 549 198 619
rect -685 516 -674 549
rect -307 516 -180 549
rect 187 516 198 549
rect 22 511 67 516
rect -824 113 -814 508
rect -1468 103 -814 113
rect -770 449 -748 472
rect -716 449 -260 472
rect -770 116 -749 449
rect -334 116 -260 449
rect -770 100 -748 116
rect -716 100 -260 116
rect -222 100 234 472
rect 266 100 280 472
rect -679 52 -292 56
rect -679 12 -669 52
rect -302 12 -292 52
rect -192 53 198 56
rect -192 13 -180 53
rect 187 13 198 53
rect 324 29 334 692
rect 366 71 376 692
rect 1764 167 1770 2268
rect 463 165 556 167
rect 463 125 473 165
rect 547 125 556 165
rect 463 115 556 125
rect 623 157 876 167
rect 623 125 634 157
rect 706 125 794 157
rect 866 125 876 157
rect 623 115 876 125
rect 943 157 1196 167
rect 943 125 954 157
rect 1026 125 1114 157
rect 1186 125 1196 157
rect 943 115 1196 125
rect 1263 157 1516 167
rect 1263 125 1274 157
rect 1346 125 1434 157
rect 1506 125 1516 157
rect 1263 115 1516 125
rect 1583 157 1770 167
rect 1583 125 1594 157
rect 1666 125 1770 157
rect 1583 71 1770 125
rect 366 65 1770 71
rect 366 61 648 65
rect 1724 61 1770 65
rect 1810 34 1816 2268
rect 1806 29 1816 34
rect 324 25 648 29
rect 1724 25 1816 29
rect 324 19 1816 25
rect -192 12 198 13
rect -679 11 -292 12
<< via1 >>
rect -1152 1426 -1143 2365
rect -1143 1426 -1112 2365
rect -965 2324 -620 2353
rect -1053 2210 -1041 2282
rect -1041 2210 -1013 2282
rect -1053 2206 -1013 2210
rect -965 2168 -620 2324
rect -965 2136 -620 2168
rect -965 1987 -620 2136
rect -1050 1906 -1010 1908
rect -1050 1836 -1041 1906
rect -1041 1836 -1010 1906
rect -1055 1718 -1015 1721
rect -1055 1646 -1041 1718
rect -1041 1646 -1015 1718
rect -1055 1645 -1015 1646
rect -375 2340 -155 2341
rect -482 2324 -155 2340
rect -482 2182 -155 2324
rect -87 2282 -47 2284
rect -87 2210 -57 2282
rect -57 2210 -47 2282
rect -87 2208 -47 2210
rect -482 2168 -320 2182
rect -482 2136 -320 2168
rect -482 1986 -320 2136
rect -88 2022 -57 2094
rect -57 2022 -48 2094
rect -475 1760 -143 1769
rect -475 1604 -143 1760
rect -88 1646 -57 1718
rect -57 1646 -48 1718
rect -475 1588 -143 1604
rect -1152 1425 -1112 1426
rect 413 2365 1798 2373
rect -509 1306 -296 1346
rect -91 1306 -51 1346
rect -1430 721 -1359 873
rect -1293 768 -1253 875
rect -1105 661 -1023 974
rect -179 1149 188 1157
rect -179 1117 187 1149
rect 187 1117 188 1149
rect -1292 384 -1232 429
rect -1232 384 -1202 429
rect -1310 307 -1306 329
rect -1306 307 -1274 329
rect -1274 307 -1270 329
rect -1310 257 -1270 307
rect -748 713 -716 1046
rect -716 713 -333 1046
rect 331 692 334 2364
rect 334 2333 371 2364
rect 413 2333 1798 2365
rect 334 692 366 2333
rect 366 692 371 2333
rect 413 2325 1774 2333
rect 1774 2325 1798 2333
rect 31 619 184 643
rect 31 549 184 619
rect 31 521 184 549
rect -749 116 -748 449
rect -748 116 -716 449
rect -716 116 -334 449
rect -669 19 -302 52
rect -669 12 -302 19
rect -180 52 187 53
rect -180 19 187 52
rect -180 13 187 19
rect 473 157 547 165
rect 473 125 474 157
rect 474 125 546 157
rect 546 125 547 157
rect 648 61 1724 65
rect 1770 61 1774 2268
rect 1774 61 1806 2268
rect 648 29 1724 61
rect 1770 34 1806 61
rect 1806 34 1810 2268
rect 648 25 1724 29
<< metal2 >>
rect -1161 2365 -1103 2378
rect 620 2373 1816 2374
rect -1161 1425 -1152 2365
rect -1112 1425 -1103 2365
rect -965 2353 -129 2370
rect -1053 2282 -1008 2320
rect -1013 2206 -1008 2282
rect -1053 2165 -1008 2206
rect -620 2341 -129 2353
rect -620 2340 -375 2341
rect -620 1987 -482 2340
rect -155 2182 -129 2341
rect 322 2364 413 2373
rect -965 1986 -482 1987
rect -320 2148 -129 2182
rect -87 2284 -5 2323
rect -47 2208 -5 2284
rect -87 2145 -5 2208
rect -965 1977 -320 1986
rect -273 2094 -48 2103
rect -273 2022 -88 2094
rect -273 2012 -48 2022
rect -965 1976 -620 1977
rect -273 1919 -182 2012
rect -1061 1908 -182 1919
rect -1061 1836 -1050 1908
rect -1010 1836 -182 1908
rect -1061 1828 -182 1836
rect -1059 1721 -999 1771
rect -1059 1645 -1055 1721
rect -1015 1645 -999 1721
rect -1059 1603 -999 1645
rect -1161 1412 -1103 1425
rect -772 1136 -562 1828
rect -486 1769 -133 1779
rect -486 1588 -475 1769
rect -143 1588 -133 1769
rect -91 1718 -48 1728
rect -91 1646 -88 1718
rect -91 1632 -48 1646
rect -486 1580 -139 1588
rect -228 1579 -139 1580
rect -512 1390 -293 1400
rect -512 1346 -501 1390
rect -302 1346 -293 1390
rect -512 1306 -509 1346
rect -296 1306 -293 1346
rect -512 1218 -501 1306
rect -302 1218 -293 1306
rect -512 1208 -293 1218
rect -223 1166 -139 1579
rect -91 1346 -51 1632
rect -91 1297 -51 1306
rect -223 1164 -32 1166
rect -223 1157 198 1164
rect -473 1136 -298 1141
rect -773 1113 -298 1136
rect -1406 1061 -298 1113
rect -1406 883 -1354 1061
rect -771 1046 -298 1061
rect -1115 974 -1013 984
rect -1440 873 -1349 883
rect -1440 721 -1430 873
rect -1359 721 -1349 873
rect -1440 711 -1349 721
rect -1303 875 -1242 885
rect -1303 768 -1293 875
rect -1253 768 -1242 875
rect -1303 440 -1242 768
rect -1115 661 -1105 974
rect -1023 661 -1013 974
rect -1115 651 -1013 661
rect -771 713 -748 1046
rect -333 713 -298 1046
rect -771 449 -298 713
rect -1303 429 -1186 440
rect -1303 384 -1292 429
rect -1202 384 -1186 429
rect -1303 372 -1186 384
rect -1322 329 -1259 330
rect -1322 257 -1310 329
rect -1270 294 -1259 329
rect -1270 257 -932 294
rect -1322 226 -932 257
rect -1000 52 -932 226
rect -771 116 -749 449
rect -334 116 -298 449
rect -771 108 -298 116
rect -223 1117 -179 1157
rect 188 1117 198 1157
rect -223 1100 198 1117
rect -223 695 196 1100
rect -223 443 -20 695
rect 322 692 331 2364
rect 371 2325 413 2364
rect 1798 2325 1816 2373
rect 371 2268 1816 2325
rect 371 692 1770 2268
rect 22 643 194 653
rect 22 521 31 643
rect 184 614 194 643
rect 460 614 556 616
rect 184 521 556 614
rect 22 518 556 521
rect 22 511 194 518
rect -223 56 198 443
rect 460 165 556 518
rect 460 125 473 165
rect 547 125 556 165
rect 460 116 556 125
rect 620 340 1770 692
rect -681 53 198 56
rect -681 52 -180 53
rect -1000 12 -669 52
rect -302 13 -180 52
rect 187 13 198 53
rect 620 105 915 340
rect 1529 105 1770 340
rect 620 65 1770 105
rect 620 25 648 65
rect 1724 34 1770 65
rect 1810 34 1816 2268
rect 1724 25 1816 34
rect 620 19 1816 25
rect -302 12 198 13
rect -681 11 198 12
<< via2 >>
rect -501 1346 -302 1390
rect -501 1306 -302 1346
rect -501 1218 -302 1306
rect 915 105 1529 340
<< metal3 >>
rect -802 1654 -294 1680
rect -802 1291 -788 1654
rect -431 1400 -294 1654
rect -431 1390 -293 1400
rect -802 1280 -501 1291
rect -512 1218 -501 1280
rect -302 1218 -293 1390
rect -512 1208 -293 1218
rect 898 340 1553 359
rect 898 105 915 340
rect 1529 105 1553 340
rect 898 93 1553 105
<< via3 >>
rect -788 1390 -431 1654
rect -788 1291 -501 1390
rect -501 1291 -431 1390
rect 915 105 1529 340
<< metal4 >>
rect -828 1654 -397 1686
rect -828 1291 -788 1654
rect -431 1291 -397 1654
rect -828 1268 -397 1291
rect 898 340 1553 359
rect 898 105 915 340
rect 1529 105 1553 340
rect 898 93 1553 105
<< via4 >>
rect -782 1300 -443 1640
rect 915 105 1529 340
<< metal5 >>
rect -814 1640 -398 1681
rect -814 1300 -782 1640
rect -443 1300 -398 1640
rect -814 1268 -398 1300
rect -69 379 1571 2019
rect 871 340 1571 379
rect 871 105 915 340
rect 1529 105 1571 340
rect 871 76 1571 105
<< via5 >>
rect -756 1311 -488 1611
<< mimcap >>
rect 51 1839 1451 1899
rect 51 559 111 1839
rect 1391 559 1451 1839
rect 51 499 1451 559
<< mimcapcontact >>
rect 111 559 1391 1839
<< metal6 >>
rect 99 1839 1403 1851
rect -89 1730 111 1839
rect -814 1683 111 1730
rect -838 1611 111 1683
rect -838 1311 -756 1611
rect -488 1311 111 1611
rect -838 1273 111 1311
rect -838 1244 -418 1273
rect -89 559 111 1273
rect 1391 559 1403 1839
rect 99 547 1403 559
<< labels >>
flabel metal2 -1157 1415 -1105 2375 1 FreeSans 320 0 0 0 VCC
port 0 n power default
flabel metal2 733 46 1782 2346 0 FreeSans 320 0 0 0 GND
port 1 nsew power default
flabel metal2 -1059 1603 -999 1771 0 FreeSans 320 0 0 0 Ibias_1u_1
port 6 nsew
flabel metal2 -1053 2165 -1008 2320 0 FreeSans 320 0 0 0 Ibias_1u_2
port 7 nsew
flabel metal2 -87 2145 -5 2323 0 FreeSans 320 0 0 0 Ibias_1u_3
port 8 nsew
flabel metal2 -1115 651 -1013 984 0 FreeSans 320 0 0 0 por
port 9 nsew
<< end >>
