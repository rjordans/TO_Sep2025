magic
tech ihp-sg13g2
magscale 1 2
timestamp 1756729118
<< nwell >>
rect 608 1566 1570 2016
rect 608 996 2682 1566
rect -1658 -8 2682 996
<< hvnmos >>
rect -1416 2468 -1216 2868
rect -1032 2468 -832 2868
rect -648 2468 -448 2868
rect -264 2468 -64 2868
rect 120 2468 320 2868
rect -1416 1890 -1216 2290
rect -1032 1890 -832 2290
rect -648 1890 -448 2290
rect -264 1890 -64 2290
rect 120 1890 320 2290
rect -1416 1312 -1216 1712
rect -1032 1312 -832 1712
rect -648 1312 -448 1712
rect -264 1312 -64 1712
rect 120 1312 320 1712
rect 896 2308 986 2368
rect 1172 2308 1262 2368
<< hvpmos >>
rect 914 1670 994 1730
rect 1172 1670 1252 1730
rect -1380 298 -1180 698
rect -1092 298 -892 698
rect -804 298 -604 698
rect -516 298 -316 698
rect -228 298 -28 698
rect 60 298 260 698
rect 902 278 982 1278
rect 1058 278 1138 1278
rect 1214 278 1294 1278
rect 1370 278 1450 1278
rect 1526 278 1606 1278
rect 1682 278 1762 1278
rect 1838 278 1918 1278
rect 1994 278 2074 1278
rect 2150 278 2230 1278
rect 2306 278 2386 1278
<< hvndiff >>
rect -1416 2922 -1216 2936
rect -1416 2890 -1402 2922
rect -1230 2890 -1216 2922
rect -1416 2868 -1216 2890
rect -1032 2922 -832 2936
rect -1032 2890 -1018 2922
rect -846 2890 -832 2922
rect -1032 2868 -832 2890
rect -648 2922 -448 2936
rect -648 2890 -634 2922
rect -462 2890 -448 2922
rect -648 2868 -448 2890
rect -264 2922 -64 2936
rect -264 2890 -250 2922
rect -78 2890 -64 2922
rect -264 2868 -64 2890
rect 120 2922 320 2936
rect 120 2890 134 2922
rect 306 2890 320 2922
rect 120 2868 320 2890
rect -1416 2446 -1216 2468
rect -1416 2414 -1402 2446
rect -1230 2414 -1216 2446
rect -1416 2400 -1216 2414
rect -1032 2446 -832 2468
rect -1032 2414 -1018 2446
rect -846 2414 -832 2446
rect -1032 2400 -832 2414
rect -648 2446 -448 2468
rect -648 2414 -634 2446
rect -462 2414 -448 2446
rect -648 2400 -448 2414
rect -264 2446 -64 2468
rect -264 2414 -250 2446
rect -78 2414 -64 2446
rect -264 2400 -64 2414
rect 120 2446 320 2468
rect 120 2414 134 2446
rect 306 2414 320 2446
rect 120 2400 320 2414
rect -1416 2344 -1216 2358
rect -1416 2312 -1402 2344
rect -1230 2312 -1216 2344
rect -1416 2290 -1216 2312
rect -1032 2344 -832 2358
rect -1032 2312 -1018 2344
rect -846 2312 -832 2344
rect -1032 2290 -832 2312
rect -648 2344 -448 2358
rect -648 2312 -634 2344
rect -462 2312 -448 2344
rect -648 2290 -448 2312
rect -264 2344 -64 2358
rect -264 2312 -250 2344
rect -78 2312 -64 2344
rect -264 2290 -64 2312
rect 120 2344 320 2358
rect 120 2312 134 2344
rect 306 2312 320 2344
rect 120 2290 320 2312
rect -1416 1868 -1216 1890
rect -1416 1836 -1402 1868
rect -1230 1836 -1216 1868
rect -1416 1822 -1216 1836
rect -1032 1868 -832 1890
rect -1032 1836 -1018 1868
rect -846 1836 -832 1868
rect -1032 1822 -832 1836
rect -648 1868 -448 1890
rect -648 1836 -634 1868
rect -462 1836 -448 1868
rect -648 1822 -448 1836
rect -264 1868 -64 1890
rect -264 1836 -250 1868
rect -78 1836 -64 1868
rect -264 1822 -64 1836
rect 120 1868 320 1890
rect 120 1836 134 1868
rect 306 1836 320 1868
rect 120 1822 320 1836
rect -1416 1766 -1216 1780
rect -1416 1734 -1402 1766
rect -1230 1734 -1216 1766
rect -1416 1712 -1216 1734
rect -1032 1766 -832 1780
rect -1032 1734 -1018 1766
rect -846 1734 -832 1766
rect -1032 1712 -832 1734
rect -648 1766 -448 1780
rect -648 1734 -634 1766
rect -462 1734 -448 1766
rect -648 1712 -448 1734
rect -264 1766 -64 1780
rect -264 1734 -250 1766
rect -78 1734 -64 1766
rect -264 1712 -64 1734
rect 120 1766 320 1780
rect 120 1734 134 1766
rect 306 1734 320 1766
rect 120 1712 320 1734
rect -1416 1290 -1216 1312
rect -1416 1258 -1402 1290
rect -1230 1258 -1216 1290
rect -1416 1244 -1216 1258
rect -1032 1290 -832 1312
rect -1032 1258 -1018 1290
rect -846 1258 -832 1290
rect -1032 1244 -832 1258
rect -648 1290 -448 1312
rect -648 1258 -634 1290
rect -462 1258 -448 1290
rect -648 1244 -448 1258
rect -264 1290 -64 1312
rect -264 1258 -250 1290
rect -78 1258 -64 1290
rect -264 1244 -64 1258
rect 120 1290 320 1312
rect 120 1258 134 1290
rect 306 1258 320 1290
rect 120 1244 320 1258
rect 828 2354 896 2368
rect 828 2322 842 2354
rect 874 2322 896 2354
rect 828 2308 896 2322
rect 986 2354 1172 2368
rect 986 2322 1008 2354
rect 1150 2322 1172 2354
rect 986 2308 1172 2322
rect 1262 2354 1330 2368
rect 1262 2322 1284 2354
rect 1316 2322 1330 2354
rect 1262 2308 1330 2322
<< hvpdiff >>
rect 846 1716 914 1730
rect 846 1684 860 1716
rect 892 1684 914 1716
rect 846 1670 914 1684
rect 994 1716 1172 1730
rect 994 1684 1020 1716
rect 1150 1684 1172 1716
rect 994 1670 1172 1684
rect 1252 1716 1332 1730
rect 1252 1684 1286 1716
rect 1318 1684 1332 1716
rect 1252 1670 1332 1684
rect -1380 752 -1180 770
rect -1380 720 -1366 752
rect -1194 720 -1180 752
rect -1380 698 -1180 720
rect -1092 752 -892 770
rect -1092 720 -1078 752
rect -906 720 -892 752
rect -1092 698 -892 720
rect -804 752 -604 770
rect -804 720 -790 752
rect -618 720 -604 752
rect -804 698 -604 720
rect -516 752 -316 770
rect -516 720 -502 752
rect -330 720 -316 752
rect -516 698 -316 720
rect -228 752 -28 770
rect -228 720 -214 752
rect -42 720 -28 752
rect -228 698 -28 720
rect 60 752 260 770
rect 60 720 74 752
rect 246 720 260 752
rect 60 698 260 720
rect -1380 266 -1180 298
rect -1380 234 -1366 266
rect -1194 234 -1180 266
rect -1380 220 -1180 234
rect -1092 266 -892 298
rect -1092 234 -1078 266
rect -906 234 -892 266
rect -1092 220 -892 234
rect -804 266 -604 298
rect -804 234 -790 266
rect -618 234 -604 266
rect -804 220 -604 234
rect -516 266 -316 298
rect -516 234 -502 266
rect -330 234 -316 266
rect -516 220 -316 234
rect -228 266 -28 298
rect -228 234 -214 266
rect -42 234 -28 266
rect -228 220 -28 234
rect 60 268 260 298
rect 60 236 74 268
rect 246 236 260 268
rect 60 222 260 236
rect 834 1254 902 1278
rect 834 298 848 1254
rect 880 298 902 1254
rect 834 278 902 298
rect 982 1256 1058 1278
rect 982 300 1004 1256
rect 1036 300 1058 1256
rect 982 278 1058 300
rect 1138 1256 1214 1278
rect 1138 300 1160 1256
rect 1192 300 1214 1256
rect 1138 278 1214 300
rect 1294 1256 1370 1278
rect 1294 300 1316 1256
rect 1348 300 1370 1256
rect 1294 278 1370 300
rect 1450 1256 1526 1278
rect 1450 300 1472 1256
rect 1504 300 1526 1256
rect 1450 278 1526 300
rect 1606 1256 1682 1278
rect 1606 300 1628 1256
rect 1660 300 1682 1256
rect 1606 278 1682 300
rect 1762 1256 1838 1278
rect 1762 300 1784 1256
rect 1816 300 1838 1256
rect 1762 278 1838 300
rect 1918 1256 1994 1278
rect 1918 300 1940 1256
rect 1972 300 1994 1256
rect 1918 278 1994 300
rect 2074 1256 2150 1278
rect 2074 300 2096 1256
rect 2128 300 2150 1256
rect 2074 278 2150 300
rect 2230 1256 2306 1278
rect 2230 300 2252 1256
rect 2284 300 2306 1256
rect 2230 278 2306 300
rect 2386 1256 2454 1278
rect 2386 300 2408 1256
rect 2440 300 2454 1256
rect 2386 278 2454 300
<< hvndiffc >>
rect -1402 2890 -1230 2922
rect -1018 2890 -846 2922
rect -634 2890 -462 2922
rect -250 2890 -78 2922
rect 134 2890 306 2922
rect -1402 2414 -1230 2446
rect -1018 2414 -846 2446
rect -634 2414 -462 2446
rect -250 2414 -78 2446
rect 134 2414 306 2446
rect -1402 2312 -1230 2344
rect -1018 2312 -846 2344
rect -634 2312 -462 2344
rect -250 2312 -78 2344
rect 134 2312 306 2344
rect -1402 1836 -1230 1868
rect -1018 1836 -846 1868
rect -634 1836 -462 1868
rect -250 1836 -78 1868
rect 134 1836 306 1868
rect -1402 1734 -1230 1766
rect -1018 1734 -846 1766
rect -634 1734 -462 1766
rect -250 1734 -78 1766
rect 134 1734 306 1766
rect -1402 1258 -1230 1290
rect -1018 1258 -846 1290
rect -634 1258 -462 1290
rect -250 1258 -78 1290
rect 134 1258 306 1290
rect 842 2322 874 2354
rect 1008 2322 1150 2354
rect 1284 2322 1316 2354
<< hvpdiffc >>
rect 860 1684 892 1716
rect 1020 1684 1150 1716
rect 1286 1684 1318 1716
rect -1366 720 -1194 752
rect -1078 720 -906 752
rect -790 720 -618 752
rect -502 720 -330 752
rect -214 720 -42 752
rect 74 720 246 752
rect -1366 234 -1194 266
rect -1078 234 -906 266
rect -790 234 -618 266
rect -502 234 -330 266
rect -214 234 -42 266
rect 74 236 246 268
rect 848 298 880 1254
rect 1004 300 1036 1256
rect 1160 300 1192 1256
rect 1316 300 1348 1256
rect 1472 300 1504 1256
rect 1628 300 1660 1256
rect 1784 300 1816 1256
rect 1940 300 1972 1256
rect 2096 300 2128 1256
rect 2252 300 2284 1256
rect 2408 300 2440 1256
<< psubdiff >>
rect -1698 -85 2682 -71
rect -1698 -1214 -1684 -85
rect -1652 -131 2636 -117
rect -1652 -1168 -1638 -131
rect 2622 -1168 2636 -131
rect -1652 -1182 2636 -1168
rect 2668 -1214 2682 -85
rect -1698 -1228 2682 -1214
<< hvpsubdiff >>
rect -1602 3026 480 3040
rect -1602 1152 -1588 3026
rect -1556 2980 434 2994
rect -1556 1198 -1542 2980
rect 420 1198 434 2980
rect -1556 1184 434 1198
rect 466 1152 480 3026
rect 726 2526 1432 2540
rect 726 2154 740 2526
rect 772 2480 1386 2494
rect 772 2200 786 2480
rect 1372 2200 1386 2480
rect 772 2186 1386 2200
rect 1418 2154 1432 2526
rect 726 2140 1432 2154
rect -1602 1138 480 1152
<< hvnsubdiff >>
rect 744 1878 1434 1892
rect 744 1522 758 1878
rect 790 1832 1388 1846
rect 790 1568 804 1832
rect 1374 1568 1388 1832
rect 790 1554 1388 1568
rect 1420 1522 1434 1878
rect 744 1508 1434 1522
rect 732 1428 2558 1442
rect -1534 858 426 872
rect -1534 130 -1520 858
rect -1488 812 380 826
rect -1488 176 -1466 812
rect 358 176 380 812
rect -1488 162 380 176
rect 412 130 426 858
rect -1534 116 426 130
rect 732 130 746 1428
rect 778 1382 2512 1396
rect 778 176 792 1382
rect 2498 176 2512 1382
rect 778 162 2512 176
rect 2544 130 2558 1428
rect 732 116 2558 130
<< psubdiffcont >>
rect -1684 -117 2668 -85
rect -1684 -1182 -1652 -117
rect 2636 -1182 2668 -117
rect -1684 -1214 2668 -1182
<< hvpsubdiffcont >>
rect -1588 2994 466 3026
rect -1588 1184 -1556 2994
rect 434 1184 466 2994
rect -1588 1152 466 1184
rect 740 2494 1418 2526
rect 740 2186 772 2494
rect 1386 2186 1418 2494
rect 740 2154 1418 2186
<< hvnsubdiffcont >>
rect 758 1846 1420 1878
rect 758 1554 790 1846
rect 1388 1554 1420 1846
rect 758 1522 1420 1554
rect -1520 826 412 858
rect -1520 162 -1488 826
rect 380 162 412 826
rect -1520 130 412 162
rect 746 1396 2544 1428
rect 746 162 778 1396
rect 2512 162 2544 1396
rect 746 130 2544 162
<< poly >>
rect -1490 2844 -1416 2868
rect -1490 2482 -1476 2844
rect -1444 2482 -1416 2844
rect -1490 2468 -1416 2482
rect -1216 2844 -1142 2868
rect -1216 2482 -1188 2844
rect -1156 2482 -1142 2844
rect -1216 2468 -1142 2482
rect -1106 2834 -1032 2868
rect -1106 2502 -1092 2834
rect -1060 2502 -1032 2834
rect -1106 2468 -1032 2502
rect -832 2834 -758 2868
rect -832 2502 -804 2834
rect -772 2502 -758 2834
rect -832 2468 -758 2502
rect -722 2834 -648 2868
rect -722 2502 -708 2834
rect -676 2502 -648 2834
rect -722 2468 -648 2502
rect -448 2834 -374 2868
rect -448 2502 -420 2834
rect -388 2502 -374 2834
rect -448 2468 -374 2502
rect -338 2834 -264 2868
rect -338 2502 -324 2834
rect -292 2502 -264 2834
rect -338 2468 -264 2502
rect -64 2834 10 2868
rect -64 2502 -36 2834
rect -4 2502 10 2834
rect -64 2468 10 2502
rect 46 2844 120 2868
rect 46 2482 60 2844
rect 92 2482 120 2844
rect 46 2468 120 2482
rect 320 2844 394 2868
rect 320 2482 348 2844
rect 380 2482 394 2844
rect 320 2468 394 2482
rect -1490 2266 -1416 2290
rect -1490 1904 -1476 2266
rect -1444 1904 -1416 2266
rect -1490 1890 -1416 1904
rect -1216 2266 -1142 2290
rect -1216 1904 -1188 2266
rect -1156 1904 -1142 2266
rect -1216 1890 -1142 1904
rect -1106 2266 -1032 2290
rect -1106 2112 -1092 2266
rect -1060 2112 -1032 2266
rect -1106 1890 -1032 2112
rect -832 2266 -758 2290
rect -832 2112 -804 2266
rect -772 2112 -758 2266
rect -832 1890 -758 2112
rect -722 2068 -648 2290
rect -722 1914 -708 2068
rect -676 1914 -648 2068
rect -722 1890 -648 1914
rect -448 2068 -374 2290
rect -448 1914 -420 2068
rect -388 1914 -374 2068
rect -448 1890 -374 1914
rect -338 2266 -264 2290
rect -338 1924 -324 2266
rect -292 1924 -264 2266
rect -338 1890 -264 1924
rect -64 2266 10 2290
rect -64 1904 -36 2266
rect -4 1904 10 2266
rect -64 1890 10 1904
rect 46 2266 120 2290
rect 46 1904 60 2266
rect 92 1904 120 2266
rect 46 1890 120 1904
rect 320 2276 394 2290
rect 320 1904 348 2276
rect 380 1904 394 2276
rect 320 1890 394 1904
rect -1490 1698 -1416 1712
rect -1490 1336 -1476 1698
rect -1444 1336 -1416 1698
rect -1490 1312 -1416 1336
rect -1216 1698 -1142 1712
rect -1216 1336 -1188 1698
rect -1156 1336 -1142 1698
rect -1216 1312 -1142 1336
rect -1106 1698 -1032 1712
rect -1106 1336 -1092 1698
rect -1060 1336 -1032 1698
rect -1106 1312 -1032 1336
rect -832 1678 -758 1712
rect -832 1336 -804 1678
rect -772 1336 -758 1678
rect -832 1312 -758 1336
rect -722 1688 -648 1712
rect -722 1534 -708 1688
rect -676 1534 -648 1688
rect -722 1312 -648 1534
rect -448 1688 -374 1712
rect -448 1534 -420 1688
rect -388 1534 -374 1688
rect -448 1312 -374 1534
rect -338 1490 -264 1712
rect -338 1336 -324 1490
rect -292 1336 -264 1490
rect -338 1312 -264 1336
rect -64 1490 10 1712
rect -64 1336 -36 1490
rect -4 1336 10 1490
rect -64 1312 10 1336
rect 46 1698 120 1712
rect 46 1336 60 1698
rect 92 1336 120 1698
rect 46 1312 120 1336
rect 320 1698 394 1712
rect 320 1326 348 1698
rect 380 1326 394 1698
rect 320 1312 394 1326
rect 896 2428 986 2442
rect 896 2396 928 2428
rect 960 2396 986 2428
rect 896 2368 986 2396
rect 1172 2428 1262 2442
rect 1172 2396 1204 2428
rect 1236 2396 1262 2428
rect 1172 2368 1262 2396
rect 896 2278 986 2308
rect 896 2246 928 2278
rect 960 2246 986 2278
rect 896 2230 986 2246
rect 1172 2276 1262 2308
rect 1172 2244 1204 2276
rect 1236 2244 1262 2276
rect 1172 2230 1262 2244
rect 914 1790 994 1804
rect 914 1758 940 1790
rect 972 1758 994 1790
rect 914 1730 994 1758
rect 1172 1790 1252 1804
rect 1172 1758 1198 1790
rect 1230 1758 1252 1790
rect 1172 1730 1252 1758
rect 914 1642 994 1670
rect 914 1610 940 1642
rect 972 1610 994 1642
rect 914 1596 994 1610
rect 1172 1642 1252 1670
rect 1172 1610 1198 1642
rect 1230 1610 1252 1642
rect 1172 1596 1252 1610
rect -1426 298 -1380 698
rect -1180 676 -1092 698
rect -1180 316 -1152 676
rect -1120 316 -1092 676
rect -1180 298 -1092 316
rect -892 676 -804 698
rect -892 316 -864 676
rect -832 316 -804 676
rect -892 298 -804 316
rect -604 676 -516 698
rect -604 316 -576 676
rect -544 316 -516 676
rect -604 298 -516 316
rect -316 676 -228 698
rect -316 316 -288 676
rect -256 316 -228 676
rect -316 298 -228 316
rect -28 676 60 698
rect -28 316 0 676
rect 32 316 60 676
rect -28 298 60 316
rect 260 298 306 698
rect 902 1338 982 1362
rect 902 1306 926 1338
rect 958 1306 982 1338
rect 902 1278 982 1306
rect 1058 1338 1138 1362
rect 1058 1306 1082 1338
rect 1114 1306 1138 1338
rect 1058 1278 1138 1306
rect 1214 1338 1294 1362
rect 1214 1306 1238 1338
rect 1270 1306 1294 1338
rect 1214 1278 1294 1306
rect 1370 1338 1450 1362
rect 1370 1306 1394 1338
rect 1426 1306 1450 1338
rect 1370 1278 1450 1306
rect 1526 1338 1606 1362
rect 1526 1306 1550 1338
rect 1582 1306 1606 1338
rect 1526 1278 1606 1306
rect 1682 1338 1762 1362
rect 1682 1306 1706 1338
rect 1738 1306 1762 1338
rect 1682 1278 1762 1306
rect 1838 1338 1918 1362
rect 1838 1306 1862 1338
rect 1894 1306 1918 1338
rect 1838 1278 1918 1306
rect 1994 1338 2074 1362
rect 1994 1306 2018 1338
rect 2050 1306 2074 1338
rect 1994 1278 2074 1306
rect 2150 1338 2230 1362
rect 2150 1306 2174 1338
rect 2206 1306 2230 1338
rect 2150 1278 2230 1306
rect 2306 1338 2386 1362
rect 2306 1306 2330 1338
rect 2362 1306 2386 1338
rect 2306 1278 2386 1306
rect 902 250 982 278
rect 902 218 926 250
rect 958 218 982 250
rect 902 204 982 218
rect 1058 250 1138 278
rect 1058 218 1082 250
rect 1114 218 1138 250
rect 1058 204 1138 218
rect 1214 250 1294 278
rect 1214 218 1238 250
rect 1270 218 1294 250
rect 1214 204 1294 218
rect 1370 250 1450 278
rect 1370 218 1394 250
rect 1426 218 1450 250
rect 1370 204 1450 218
rect 1526 250 1606 278
rect 1526 218 1550 250
rect 1582 218 1606 250
rect 1526 204 1606 218
rect 1682 250 1762 278
rect 1682 218 1706 250
rect 1738 218 1762 250
rect 1682 204 1762 218
rect 1838 250 1918 278
rect 1838 218 1862 250
rect 1894 218 1918 250
rect 1838 204 1918 218
rect 1994 250 2074 278
rect 1994 218 2018 250
rect 2050 218 2074 250
rect 1994 204 2074 218
rect 2150 250 2230 278
rect 2150 218 2174 250
rect 2206 218 2230 250
rect 2150 204 2230 218
rect 2306 250 2386 278
rect 2306 218 2330 250
rect 2362 218 2386 250
rect 2306 204 2386 218
rect -1558 -178 -1458 -164
rect -1558 -210 -1544 -178
rect -1472 -210 -1458 -178
rect -1558 -250 -1458 -210
rect -1558 -1090 -1458 -1050
rect -1558 -1122 -1544 -1090
rect -1472 -1122 -1458 -1090
rect -1558 -1136 -1458 -1122
rect -1398 -178 -1298 -164
rect -1398 -210 -1384 -178
rect -1312 -210 -1298 -178
rect -1398 -250 -1298 -210
rect -1398 -1090 -1298 -1050
rect -1398 -1122 -1384 -1090
rect -1312 -1122 -1298 -1090
rect -1398 -1136 -1298 -1122
rect -1238 -178 -1138 -164
rect -1238 -210 -1224 -178
rect -1152 -210 -1138 -178
rect -1238 -250 -1138 -210
rect -1238 -1090 -1138 -1050
rect -1238 -1122 -1224 -1090
rect -1152 -1122 -1138 -1090
rect -1238 -1136 -1138 -1122
rect -1078 -178 -978 -164
rect -1078 -210 -1064 -178
rect -992 -210 -978 -178
rect -1078 -250 -978 -210
rect -1078 -1090 -978 -1050
rect -1078 -1122 -1064 -1090
rect -992 -1122 -978 -1090
rect -1078 -1136 -978 -1122
rect -918 -178 -818 -164
rect -918 -210 -904 -178
rect -832 -210 -818 -178
rect -918 -250 -818 -210
rect -918 -1090 -818 -1050
rect -918 -1122 -904 -1090
rect -832 -1122 -818 -1090
rect -918 -1136 -818 -1122
rect -758 -178 -658 -164
rect -758 -210 -744 -178
rect -672 -210 -658 -178
rect -758 -250 -658 -210
rect -758 -1090 -658 -1050
rect -758 -1122 -744 -1090
rect -672 -1122 -658 -1090
rect -758 -1136 -658 -1122
rect -598 -178 -498 -164
rect -598 -210 -584 -178
rect -512 -210 -498 -178
rect -598 -250 -498 -210
rect -598 -1090 -498 -1050
rect -598 -1122 -584 -1090
rect -512 -1122 -498 -1090
rect -598 -1136 -498 -1122
rect -438 -178 -338 -164
rect -438 -210 -424 -178
rect -352 -210 -338 -178
rect -438 -250 -338 -210
rect -438 -1090 -338 -1050
rect -438 -1122 -424 -1090
rect -352 -1122 -338 -1090
rect -438 -1136 -338 -1122
rect -278 -178 -178 -164
rect -278 -210 -264 -178
rect -192 -210 -178 -178
rect -278 -250 -178 -210
rect -278 -1090 -178 -1050
rect -278 -1122 -264 -1090
rect -192 -1122 -178 -1090
rect -278 -1136 -178 -1122
rect -118 -178 -18 -164
rect -118 -210 -104 -178
rect -32 -210 -18 -178
rect -118 -250 -18 -210
rect -118 -1090 -18 -1050
rect -118 -1122 -104 -1090
rect -32 -1122 -18 -1090
rect -118 -1136 -18 -1122
rect 42 -178 142 -164
rect 42 -210 56 -178
rect 128 -210 142 -178
rect 42 -250 142 -210
rect 42 -1090 142 -1050
rect 42 -1122 56 -1090
rect 128 -1122 142 -1090
rect 42 -1136 142 -1122
rect 202 -178 302 -164
rect 202 -210 216 -178
rect 288 -210 302 -178
rect 202 -250 302 -210
rect 202 -1090 302 -1050
rect 202 -1122 216 -1090
rect 288 -1122 302 -1090
rect 202 -1136 302 -1122
rect 362 -178 462 -164
rect 362 -210 376 -178
rect 448 -210 462 -178
rect 362 -250 462 -210
rect 362 -1090 462 -1050
rect 362 -1122 376 -1090
rect 448 -1122 462 -1090
rect 362 -1136 462 -1122
rect 522 -178 622 -164
rect 522 -210 536 -178
rect 608 -210 622 -178
rect 522 -250 622 -210
rect 522 -1090 622 -1050
rect 522 -1122 536 -1090
rect 608 -1122 622 -1090
rect 522 -1136 622 -1122
rect 682 -178 782 -164
rect 682 -210 696 -178
rect 768 -210 782 -178
rect 682 -250 782 -210
rect 682 -1090 782 -1050
rect 682 -1122 696 -1090
rect 768 -1122 782 -1090
rect 682 -1136 782 -1122
rect 842 -178 942 -164
rect 842 -210 856 -178
rect 928 -210 942 -178
rect 842 -250 942 -210
rect 842 -1090 942 -1050
rect 842 -1122 856 -1090
rect 928 -1122 942 -1090
rect 842 -1136 942 -1122
rect 1002 -178 1102 -164
rect 1002 -210 1016 -178
rect 1088 -210 1102 -178
rect 1002 -250 1102 -210
rect 1002 -1090 1102 -1050
rect 1002 -1122 1016 -1090
rect 1088 -1122 1102 -1090
rect 1002 -1136 1102 -1122
rect 1162 -178 1262 -164
rect 1162 -210 1176 -178
rect 1248 -210 1262 -178
rect 1162 -250 1262 -210
rect 1162 -1090 1262 -1050
rect 1162 -1122 1176 -1090
rect 1248 -1122 1262 -1090
rect 1162 -1136 1262 -1122
rect 1322 -178 1422 -164
rect 1322 -210 1336 -178
rect 1408 -210 1422 -178
rect 1322 -250 1422 -210
rect 1322 -1090 1422 -1050
rect 1322 -1122 1336 -1090
rect 1408 -1122 1422 -1090
rect 1322 -1136 1422 -1122
rect 1482 -178 1582 -164
rect 1482 -210 1496 -178
rect 1568 -210 1582 -178
rect 1482 -250 1582 -210
rect 1482 -1090 1582 -1050
rect 1482 -1122 1496 -1090
rect 1568 -1122 1582 -1090
rect 1482 -1136 1582 -1122
rect 1642 -178 1742 -164
rect 1642 -210 1656 -178
rect 1728 -210 1742 -178
rect 1642 -250 1742 -210
rect 1642 -1090 1742 -1050
rect 1642 -1122 1656 -1090
rect 1728 -1122 1742 -1090
rect 1642 -1136 1742 -1122
rect 1802 -178 1902 -164
rect 1802 -210 1816 -178
rect 1888 -210 1902 -178
rect 1802 -250 1902 -210
rect 1802 -1090 1902 -1050
rect 1802 -1122 1816 -1090
rect 1888 -1122 1902 -1090
rect 1802 -1136 1902 -1122
rect 1962 -178 2062 -164
rect 1962 -210 1976 -178
rect 2048 -210 2062 -178
rect 1962 -250 2062 -210
rect 1962 -1090 2062 -1050
rect 1962 -1122 1976 -1090
rect 2048 -1122 2062 -1090
rect 1962 -1136 2062 -1122
rect 2122 -178 2222 -164
rect 2122 -210 2136 -178
rect 2208 -210 2222 -178
rect 2122 -250 2222 -210
rect 2122 -1090 2222 -1050
rect 2122 -1122 2136 -1090
rect 2208 -1122 2222 -1090
rect 2122 -1136 2222 -1122
rect 2282 -178 2382 -164
rect 2282 -210 2296 -178
rect 2368 -210 2382 -178
rect 2282 -250 2382 -210
rect 2282 -1090 2382 -1050
rect 2282 -1122 2296 -1090
rect 2368 -1122 2382 -1090
rect 2282 -1136 2382 -1122
rect 2442 -178 2542 -164
rect 2442 -210 2456 -178
rect 2528 -210 2542 -178
rect 2442 -250 2542 -210
rect 2442 -1090 2542 -1050
rect 2442 -1122 2456 -1090
rect 2528 -1122 2542 -1090
rect 2442 -1136 2542 -1122
<< polycont >>
rect -1476 2482 -1444 2844
rect -1188 2482 -1156 2844
rect -1092 2502 -1060 2834
rect -804 2502 -772 2834
rect -708 2502 -676 2834
rect -420 2502 -388 2834
rect -324 2502 -292 2834
rect -36 2502 -4 2834
rect 60 2482 92 2844
rect 348 2482 380 2844
rect -1476 1904 -1444 2266
rect -1188 1904 -1156 2266
rect -1092 2112 -1060 2266
rect -804 2112 -772 2266
rect -708 1914 -676 2068
rect -420 1914 -388 2068
rect -324 1924 -292 2266
rect -36 1904 -4 2266
rect 60 1904 92 2266
rect 348 1904 380 2276
rect -1476 1336 -1444 1698
rect -1188 1336 -1156 1698
rect -1092 1336 -1060 1698
rect -804 1336 -772 1678
rect -708 1534 -676 1688
rect -420 1534 -388 1688
rect -324 1336 -292 1490
rect -36 1336 -4 1490
rect 60 1336 92 1698
rect 348 1326 380 1698
rect 928 2396 960 2428
rect 1204 2396 1236 2428
rect 928 2246 960 2278
rect 1204 2244 1236 2276
rect 940 1758 972 1790
rect 1198 1758 1230 1790
rect 940 1610 972 1642
rect 1198 1610 1230 1642
rect -1152 316 -1120 676
rect -864 316 -832 676
rect -576 316 -544 676
rect -288 316 -256 676
rect 0 316 32 676
rect 926 1306 958 1338
rect 1082 1306 1114 1338
rect 1238 1306 1270 1338
rect 1394 1306 1426 1338
rect 1550 1306 1582 1338
rect 1706 1306 1738 1338
rect 1862 1306 1894 1338
rect 2018 1306 2050 1338
rect 2174 1306 2206 1338
rect 2330 1306 2362 1338
rect 926 218 958 250
rect 1082 218 1114 250
rect 1238 218 1270 250
rect 1394 218 1426 250
rect 1550 218 1582 250
rect 1706 218 1738 250
rect 1862 218 1894 250
rect 2018 218 2050 250
rect 2174 218 2206 250
rect 2330 218 2362 250
rect -1544 -210 -1472 -178
rect -1544 -1122 -1472 -1090
rect -1384 -210 -1312 -178
rect -1384 -1122 -1312 -1090
rect -1224 -210 -1152 -178
rect -1224 -1122 -1152 -1090
rect -1064 -210 -992 -178
rect -1064 -1122 -992 -1090
rect -904 -210 -832 -178
rect -904 -1122 -832 -1090
rect -744 -210 -672 -178
rect -744 -1122 -672 -1090
rect -584 -210 -512 -178
rect -584 -1122 -512 -1090
rect -424 -210 -352 -178
rect -424 -1122 -352 -1090
rect -264 -210 -192 -178
rect -264 -1122 -192 -1090
rect -104 -210 -32 -178
rect -104 -1122 -32 -1090
rect 56 -210 128 -178
rect 56 -1122 128 -1090
rect 216 -210 288 -178
rect 216 -1122 288 -1090
rect 376 -210 448 -178
rect 376 -1122 448 -1090
rect 536 -210 608 -178
rect 536 -1122 608 -1090
rect 696 -210 768 -178
rect 696 -1122 768 -1090
rect 856 -210 928 -178
rect 856 -1122 928 -1090
rect 1016 -210 1088 -178
rect 1016 -1122 1088 -1090
rect 1176 -210 1248 -178
rect 1176 -1122 1248 -1090
rect 1336 -210 1408 -178
rect 1336 -1122 1408 -1090
rect 1496 -210 1568 -178
rect 1496 -1122 1568 -1090
rect 1656 -210 1728 -178
rect 1656 -1122 1728 -1090
rect 1816 -210 1888 -178
rect 1816 -1122 1888 -1090
rect 1976 -210 2048 -178
rect 1976 -1122 2048 -1090
rect 2136 -210 2208 -178
rect 2136 -1122 2208 -1090
rect 2296 -210 2368 -178
rect 2296 -1122 2368 -1090
rect 2456 -210 2528 -178
rect 2456 -1122 2528 -1090
<< xpolyres >>
rect -1558 -1050 -1458 -250
rect -1398 -1050 -1298 -250
rect -1238 -1050 -1138 -250
rect -1078 -1050 -978 -250
rect -918 -1050 -818 -250
rect -758 -1050 -658 -250
rect -598 -1050 -498 -250
rect -438 -1050 -338 -250
rect -278 -1050 -178 -250
rect -118 -1050 -18 -250
rect 42 -1050 142 -250
rect 202 -1050 302 -250
rect 362 -1050 462 -250
rect 522 -1050 622 -250
rect 682 -1050 782 -250
rect 842 -1050 942 -250
rect 1002 -1050 1102 -250
rect 1162 -1050 1262 -250
rect 1322 -1050 1422 -250
rect 1482 -1050 1582 -250
rect 1642 -1050 1742 -250
rect 1802 -1050 1902 -250
rect 1962 -1050 2062 -250
rect 2122 -1050 2222 -250
rect 2282 -1050 2382 -250
rect 2442 -1050 2542 -250
<< metal1 >>
rect -1598 3026 476 3036
rect -1598 1164 -1592 3026
rect -1552 2922 434 2994
rect -1552 2890 -1402 2922
rect -1230 2890 -1018 2922
rect -846 2890 -634 2922
rect -462 2890 -250 2922
rect -78 2890 134 2922
rect 306 2890 434 2922
rect -1552 1194 -1546 2890
rect -1402 2880 -1230 2890
rect -1018 2880 -846 2890
rect -634 2880 -462 2890
rect -250 2880 -78 2890
rect 134 2880 306 2890
rect -1476 2844 -1444 2854
rect -1476 2472 -1444 2482
rect -1400 2456 -1232 2880
rect -1188 2844 -1156 2854
rect 60 2844 92 2854
rect -1156 2834 60 2844
rect -1156 2502 -1092 2834
rect -1060 2832 -804 2834
rect -772 2832 -708 2834
rect -676 2832 -420 2834
rect -388 2832 -324 2834
rect -292 2832 -36 2834
rect -4 2832 60 2834
rect -1156 2498 -1080 2502
rect 28 2498 60 2832
rect -1156 2492 60 2498
rect -1188 2472 -1156 2482
rect -1402 2446 -1230 2456
rect -1402 2404 -1230 2414
rect -1018 2446 -846 2456
rect -1018 2354 -846 2414
rect -644 2446 -452 2492
rect 60 2472 92 2482
rect 136 2456 304 2880
rect 348 2844 380 2854
rect 348 2472 380 2482
rect -644 2414 -634 2446
rect -462 2414 -452 2446
rect -644 2404 -452 2414
rect -250 2446 -78 2456
rect -250 2354 -78 2414
rect 134 2446 306 2456
rect 134 2404 306 2414
rect -1402 2344 306 2354
rect -1230 2312 -1018 2344
rect -846 2312 -634 2344
rect -462 2312 -250 2344
rect -78 2312 134 2344
rect -1402 2302 -1230 2312
rect -1018 2302 -846 2312
rect -634 2302 -462 2312
rect -250 2302 -78 2312
rect 134 2302 306 2312
rect -1476 2266 -1444 2276
rect -1400 2256 -1232 2302
rect -1188 2266 -1156 2276
rect 60 2266 92 2276
rect -1444 1904 -1188 2256
rect -1102 2112 -1092 2266
rect -1060 2112 -804 2266
rect -772 2112 -324 2266
rect -1476 1894 -1156 1904
rect -1102 2054 -708 2068
rect -1102 1944 -1074 2054
rect -760 1944 -708 2054
rect -1102 1914 -708 1944
rect -676 1914 -420 2068
rect -388 1914 -378 2068
rect -292 2242 -36 2266
rect -292 2122 -290 2242
rect -292 1938 -98 2122
rect -292 1924 -36 1938
rect -324 1914 -36 1924
rect -1448 1868 -1180 1894
rect -1448 1836 -1402 1868
rect -1230 1836 -1180 1868
rect -1448 1766 -1180 1836
rect -1448 1734 -1402 1766
rect -1230 1734 -1180 1766
rect -1448 1708 -1180 1734
rect -1102 1708 -1064 1914
rect -4 1904 6 2266
rect -36 1894 6 1904
rect 136 2256 304 2302
rect 348 2276 380 2286
rect 92 1904 348 2256
rect 60 1894 380 1904
rect -644 1868 -454 1870
rect -250 1868 -78 1878
rect -1028 1836 -1018 1868
rect -846 1836 -728 1868
rect -1028 1826 -728 1836
rect -644 1836 -634 1868
rect -462 1836 -336 1868
rect -644 1828 -624 1836
rect -472 1828 -336 1836
rect -644 1826 -336 1828
rect -250 1828 -240 1836
rect -88 1828 -78 1836
rect -250 1826 -78 1828
rect -770 1776 -728 1826
rect -380 1776 -336 1826
rect -1018 1770 -846 1776
rect -1018 1766 -1008 1770
rect -856 1766 -846 1770
rect -770 1774 -452 1776
rect -770 1766 -628 1774
rect -476 1766 -452 1774
rect -770 1734 -634 1766
rect -462 1734 -452 1766
rect -380 1766 -68 1776
rect -380 1734 -250 1766
rect -78 1734 -68 1766
rect -1018 1730 -1008 1734
rect -856 1730 -846 1734
rect -642 1732 -452 1734
rect -1018 1724 -846 1730
rect -1476 1698 -1156 1708
rect -1444 1344 -1188 1698
rect -1476 1326 -1444 1336
rect -1400 1300 -1232 1344
rect -1102 1698 -1060 1708
rect -1102 1336 -1092 1698
rect -32 1688 6 1894
rect 80 1868 364 1894
rect 80 1836 134 1868
rect 306 1836 364 1868
rect 80 1766 364 1836
rect 80 1734 134 1766
rect 306 1734 364 1766
rect 80 1708 364 1734
rect -1060 1678 -772 1688
rect -1060 1336 -804 1678
rect -718 1534 -708 1688
rect -676 1534 -420 1688
rect -388 1534 6 1688
rect 60 1698 380 1708
rect -772 1336 -324 1490
rect -292 1336 -36 1490
rect -4 1336 6 1490
rect 92 1340 348 1698
rect -1188 1326 -1156 1336
rect 60 1326 92 1336
rect 136 1300 304 1340
rect 348 1316 380 1326
rect -1402 1290 -1230 1300
rect -1018 1290 -846 1300
rect -634 1290 -462 1300
rect -250 1290 -78 1300
rect 134 1290 306 1300
rect -1230 1258 -1018 1290
rect -846 1258 -634 1290
rect -462 1258 -250 1290
rect -78 1258 134 1290
rect -1402 1248 -1230 1258
rect -1018 1248 -846 1258
rect -634 1248 -462 1258
rect -250 1248 -78 1258
rect 134 1248 306 1258
rect 424 1194 434 2890
rect -1552 1184 434 1194
rect 466 2536 476 3026
rect 466 2526 1428 2536
rect 466 2154 740 2526
rect 772 2484 1386 2494
rect 772 2196 782 2484
rect 928 2428 960 2438
rect 832 2398 884 2410
rect 832 2358 836 2398
rect 876 2358 884 2398
rect 832 2354 884 2358
rect 832 2322 842 2354
rect 874 2322 884 2354
rect 832 2296 884 2322
rect 928 2292 960 2396
rect 1008 2354 1150 2484
rect 922 2282 966 2292
rect 922 2242 924 2282
rect 964 2242 966 2282
rect 922 2232 966 2242
rect 1008 2196 1150 2322
rect 1204 2428 1236 2438
rect 1204 2292 1236 2396
rect 1274 2358 1326 2376
rect 1274 2318 1280 2358
rect 1320 2318 1326 2358
rect 1274 2296 1326 2318
rect 1190 2282 1236 2292
rect 1190 2242 1192 2282
rect 1232 2276 1236 2282
rect 1232 2242 1236 2244
rect 1190 2232 1236 2242
rect 1376 2196 1386 2484
rect 772 2186 1386 2196
rect 1418 2154 1428 2526
rect 466 2144 1428 2154
rect -1598 1152 -1588 1164
rect 466 1152 476 2144
rect 748 1878 1430 1888
rect 748 1522 758 1878
rect 790 1836 1388 1846
rect 790 1564 800 1836
rect 940 1790 972 1800
rect 842 1762 894 1774
rect 842 1722 848 1762
rect 888 1722 894 1762
rect 842 1716 894 1722
rect 842 1684 860 1716
rect 892 1684 894 1716
rect 842 1658 894 1684
rect 940 1676 972 1758
rect 1020 1716 1150 1836
rect 1198 1790 1230 1800
rect 1190 1772 1198 1782
rect 1230 1772 1234 1782
rect 1190 1732 1192 1772
rect 1232 1732 1234 1772
rect 1190 1722 1234 1732
rect 934 1660 978 1676
rect 934 1620 936 1660
rect 976 1620 978 1660
rect 934 1610 940 1620
rect 972 1610 978 1620
rect 934 1600 978 1610
rect 1020 1564 1150 1684
rect 1198 1642 1230 1722
rect 1276 1720 1336 1742
rect 1276 1680 1282 1720
rect 1322 1680 1336 1720
rect 1276 1658 1336 1680
rect 1198 1600 1230 1610
rect 1378 1564 1388 1836
rect 790 1554 1388 1564
rect 1420 1546 1430 1878
rect 1420 1522 1432 1546
rect 748 1438 1432 1522
rect -1598 1142 476 1152
rect 736 1428 2554 1438
rect -1530 866 422 868
rect 736 866 746 1428
rect -1530 858 746 866
rect -1530 130 -1520 858
rect -1488 818 380 826
rect -1488 170 -1478 818
rect -1366 752 -1194 818
rect -1366 710 -1194 720
rect -1078 752 -906 762
rect -1078 676 -1074 720
rect -1164 316 -1152 676
rect -1120 648 -1074 676
rect -914 676 -906 720
rect -800 758 -608 762
rect -800 752 -786 758
rect -626 752 -608 758
rect -800 720 -790 752
rect -618 720 -608 752
rect -800 718 -786 720
rect -626 718 -608 720
rect -800 712 -608 718
rect -502 752 -330 762
rect -502 676 -330 720
rect -224 756 -32 762
rect -224 752 -206 756
rect -46 752 -32 756
rect -224 720 -214 752
rect -42 720 -32 752
rect -224 716 -206 720
rect -46 716 -32 720
rect -224 712 -32 716
rect 64 752 256 818
rect 64 720 74 752
rect 246 720 256 752
rect 64 712 256 720
rect -914 648 -864 676
rect -1120 316 -864 648
rect -832 316 -576 676
rect -544 316 -288 676
rect -256 316 0 676
rect 32 316 42 676
rect -1366 266 -1194 276
rect -1366 170 -1194 234
rect -1078 266 -906 276
rect -1078 170 -906 234
rect -790 266 -618 276
rect -790 170 -618 234
rect -502 266 -330 276
rect -502 170 -330 234
rect -214 266 -42 276
rect -214 170 -42 234
rect 74 268 246 278
rect 74 170 246 236
rect 370 170 380 818
rect -1488 162 380 170
rect 412 130 746 858
rect 778 1386 2512 1396
rect 778 172 788 1386
rect 848 1254 880 1386
rect 842 1242 848 1252
rect 926 1338 958 1348
rect 880 1242 886 1252
rect 842 864 844 1242
rect 884 864 886 1242
rect 842 854 848 864
rect 880 854 886 864
rect 926 816 958 1306
rect 1082 1338 1114 1348
rect 1004 1256 1036 1270
rect 920 806 964 816
rect 920 722 922 806
rect 962 722 964 806
rect 920 712 964 722
rect 848 172 880 298
rect 926 250 958 712
rect 998 664 1004 674
rect 1082 816 1114 1306
rect 1160 1256 1192 1386
rect 1154 1244 1160 1254
rect 1238 1338 1270 1348
rect 1192 1244 1198 1254
rect 1154 866 1156 1244
rect 1196 866 1198 1244
rect 1154 854 1160 866
rect 1076 806 1120 816
rect 1076 722 1078 806
rect 1118 722 1120 806
rect 1076 712 1120 722
rect 1036 664 1042 674
rect 998 286 1000 664
rect 1040 286 1042 664
rect 998 272 1042 286
rect 926 208 958 218
rect 1082 250 1114 712
rect 1082 208 1114 218
rect 1192 854 1198 866
rect 1238 816 1270 1306
rect 1394 1338 1426 1348
rect 1316 1256 1348 1270
rect 1232 806 1276 816
rect 1232 722 1234 806
rect 1274 722 1276 806
rect 1232 712 1276 722
rect 1160 172 1192 300
rect 1238 250 1270 712
rect 1310 664 1316 674
rect 1394 816 1426 1306
rect 1472 1256 1504 1386
rect 1466 1244 1472 1254
rect 1550 1338 1582 1348
rect 1504 1244 1510 1254
rect 1466 866 1468 1244
rect 1508 866 1510 1244
rect 1466 854 1472 866
rect 1388 806 1432 816
rect 1388 722 1390 806
rect 1430 722 1432 806
rect 1388 712 1432 722
rect 1348 664 1354 674
rect 1310 286 1312 664
rect 1352 286 1354 664
rect 1310 274 1354 286
rect 1238 208 1270 218
rect 1394 250 1426 712
rect 1394 208 1426 218
rect 1504 854 1510 866
rect 1550 816 1582 1306
rect 1706 1338 1738 1348
rect 1628 1256 1660 1270
rect 1544 806 1588 816
rect 1544 722 1546 806
rect 1586 722 1588 806
rect 1544 712 1588 722
rect 1472 172 1504 300
rect 1550 250 1582 712
rect 1622 664 1628 674
rect 1706 816 1738 1306
rect 1784 1256 1816 1386
rect 1778 1244 1784 1254
rect 1862 1338 1894 1348
rect 1816 1244 1822 1254
rect 1778 866 1780 1244
rect 1820 866 1822 1244
rect 1778 854 1784 866
rect 1700 806 1744 816
rect 1700 722 1702 806
rect 1742 722 1744 806
rect 1700 712 1744 722
rect 1660 664 1666 674
rect 1622 286 1624 664
rect 1664 286 1666 664
rect 1622 274 1666 286
rect 1550 208 1582 218
rect 1706 250 1738 712
rect 1706 208 1738 218
rect 1816 854 1822 866
rect 1862 816 1894 1306
rect 2018 1338 2050 1348
rect 1940 1256 1972 1270
rect 1856 806 1900 816
rect 1856 722 1858 806
rect 1898 722 1900 806
rect 1856 712 1900 722
rect 1784 172 1816 300
rect 1862 250 1894 712
rect 1934 664 1940 674
rect 2018 816 2050 1306
rect 2096 1256 2128 1386
rect 2090 1244 2096 1254
rect 2174 1338 2206 1348
rect 2128 1244 2134 1254
rect 2090 866 2092 1244
rect 2132 866 2134 1244
rect 2090 854 2096 866
rect 2012 806 2056 816
rect 2012 722 2014 806
rect 2054 722 2056 806
rect 2012 712 2056 722
rect 1972 664 1978 674
rect 1934 286 1936 664
rect 1976 286 1978 664
rect 1934 274 1978 286
rect 1862 208 1894 218
rect 2018 250 2050 712
rect 2018 208 2050 218
rect 2128 854 2134 866
rect 2174 816 2206 1306
rect 2330 1338 2362 1348
rect 2252 1256 2284 1270
rect 2168 806 2212 816
rect 2168 722 2170 806
rect 2210 722 2212 806
rect 2168 712 2212 722
rect 2096 172 2128 300
rect 2174 250 2206 712
rect 2246 664 2252 674
rect 2330 816 2362 1306
rect 2408 1256 2440 1386
rect 2402 1244 2408 1254
rect 2440 1244 2446 1254
rect 2402 866 2404 1244
rect 2444 866 2446 1244
rect 2402 852 2408 866
rect 2324 806 2368 816
rect 2324 722 2326 806
rect 2366 722 2368 806
rect 2324 712 2368 722
rect 2284 664 2290 674
rect 2246 286 2248 664
rect 2288 286 2290 664
rect 2246 274 2290 286
rect 2174 208 2206 218
rect 2330 250 2362 712
rect 2330 208 2362 218
rect 2440 852 2446 866
rect 2408 172 2440 300
rect 2502 172 2512 1386
rect 778 162 2512 172
rect 2544 130 2554 1428
rect -1530 120 2554 130
rect -1694 -85 2678 -75
rect -1694 -1214 -1684 -85
rect -1468 -127 2636 -117
rect -1468 -178 -1298 -127
rect -1468 -210 -1384 -178
rect -1312 -210 -1298 -178
rect -1468 -212 -1298 -210
rect -1652 -220 -1298 -212
rect -1238 -178 -978 -164
rect -1238 -210 -1224 -178
rect -1152 -210 -1064 -178
rect -992 -210 -978 -178
rect -1238 -220 -978 -210
rect -918 -178 -658 -164
rect -918 -210 -904 -178
rect -832 -210 -744 -178
rect -672 -210 -658 -178
rect -918 -220 -658 -210
rect -598 -178 -338 -164
rect -598 -210 -584 -178
rect -512 -210 -424 -178
rect -352 -210 -338 -178
rect -598 -220 -338 -210
rect -278 -178 -18 -164
rect -278 -210 -264 -178
rect -192 -210 -104 -178
rect -32 -210 -18 -178
rect -278 -220 -18 -210
rect 42 -178 302 -164
rect 42 -210 56 -178
rect 128 -210 216 -178
rect 288 -210 302 -178
rect 42 -220 302 -210
rect 362 -178 622 -164
rect 362 -210 376 -178
rect 448 -210 536 -178
rect 608 -210 622 -178
rect 362 -220 622 -210
rect 682 -178 942 -164
rect 682 -210 696 -178
rect 768 -210 856 -178
rect 928 -210 942 -178
rect 682 -220 942 -210
rect 1002 -178 1262 -164
rect 1002 -210 1016 -178
rect 1088 -210 1176 -178
rect 1248 -210 1262 -178
rect 1002 -220 1262 -210
rect 1322 -178 1582 -164
rect 1322 -210 1336 -178
rect 1408 -210 1496 -178
rect 1568 -210 1582 -178
rect 1322 -220 1582 -210
rect 1642 -174 1902 -164
rect 1642 -214 1656 -174
rect 1888 -214 1902 -174
rect 1642 -220 1902 -214
rect 1962 -178 2222 -164
rect 1962 -210 1976 -178
rect 2048 -210 2136 -178
rect 2208 -210 2222 -178
rect 1962 -220 2222 -210
rect 2282 -174 2382 -164
rect 2282 -214 2296 -174
rect 2368 -214 2382 -174
rect 2282 -220 2382 -214
rect 2442 -178 2636 -127
rect 2442 -210 2456 -178
rect 2528 -210 2636 -178
rect 2442 -220 2636 -210
rect -1652 -1080 -1642 -220
rect 2626 -1080 2636 -220
rect -1652 -1090 -1458 -1080
rect -1466 -1172 -1458 -1090
rect -1398 -1090 -1138 -1080
rect -1398 -1122 -1384 -1090
rect -1312 -1122 -1224 -1090
rect -1152 -1122 -1138 -1090
rect -1398 -1136 -1138 -1122
rect -1078 -1090 -818 -1080
rect -1078 -1122 -1064 -1090
rect -992 -1122 -904 -1090
rect -832 -1122 -818 -1090
rect -1078 -1136 -818 -1122
rect -758 -1090 -498 -1080
rect -758 -1122 -744 -1090
rect -672 -1122 -584 -1090
rect -512 -1122 -498 -1090
rect -758 -1136 -498 -1122
rect -438 -1090 -178 -1080
rect -438 -1122 -424 -1090
rect -352 -1122 -264 -1090
rect -192 -1122 -178 -1090
rect -438 -1136 -178 -1122
rect -118 -1090 142 -1080
rect -118 -1122 -104 -1090
rect -32 -1122 56 -1090
rect 128 -1122 142 -1090
rect -118 -1136 142 -1122
rect 202 -1090 462 -1080
rect 202 -1122 216 -1090
rect 288 -1122 376 -1090
rect 448 -1122 462 -1090
rect 202 -1136 462 -1122
rect 522 -1090 782 -1080
rect 522 -1122 536 -1090
rect 608 -1122 696 -1090
rect 768 -1122 782 -1090
rect 522 -1136 782 -1122
rect 842 -1090 1102 -1080
rect 842 -1122 856 -1090
rect 928 -1122 1016 -1090
rect 1088 -1122 1102 -1090
rect 842 -1136 1102 -1122
rect 1162 -1090 1422 -1080
rect 1162 -1122 1176 -1090
rect 1248 -1122 1336 -1090
rect 1408 -1122 1422 -1090
rect 1162 -1136 1422 -1122
rect 1482 -1090 1742 -1080
rect 1482 -1122 1496 -1090
rect 1568 -1122 1656 -1090
rect 1728 -1122 1742 -1090
rect 1482 -1136 1742 -1122
rect 1802 -1090 2062 -1080
rect 1802 -1122 1816 -1090
rect 1888 -1122 1976 -1090
rect 2048 -1122 2062 -1090
rect 1802 -1136 2062 -1122
rect 2122 -1090 2382 -1080
rect 2122 -1122 2136 -1090
rect 2208 -1122 2296 -1090
rect 2368 -1122 2382 -1090
rect 2122 -1136 2382 -1122
rect 2442 -1090 2636 -1080
rect 2442 -1122 2456 -1090
rect 2528 -1122 2636 -1090
rect 2442 -1172 2636 -1122
rect -1466 -1182 2636 -1172
rect 2668 -1214 2678 -85
rect -1694 -1224 2678 -1214
<< via1 >>
rect -1592 1164 -1588 3026
rect -1588 2994 -1552 3026
rect -1588 1184 -1556 2994
rect -1556 1184 -1552 2994
rect -1080 2502 -1060 2832
rect -1060 2502 -804 2832
rect -804 2502 -772 2832
rect -772 2502 -708 2832
rect -708 2502 -676 2832
rect -676 2502 -420 2832
rect -420 2502 -388 2832
rect -388 2502 -324 2832
rect -324 2502 -292 2832
rect -292 2502 -36 2832
rect -36 2502 -4 2832
rect -4 2502 28 2832
rect -1080 2498 28 2502
rect -1074 1944 -760 2054
rect -290 2122 -36 2242
rect -98 1938 -36 2122
rect -36 1938 -18 2242
rect -624 1836 -472 1868
rect -624 1828 -472 1836
rect -240 1836 -88 1868
rect -240 1828 -88 1836
rect -1008 1766 -856 1770
rect -1008 1734 -856 1766
rect -628 1766 -476 1774
rect -628 1734 -476 1766
rect -1008 1730 -856 1734
rect 836 2358 876 2398
rect 924 2278 964 2282
rect 924 2246 928 2278
rect 928 2246 960 2278
rect 960 2246 964 2278
rect 924 2242 964 2246
rect 1280 2354 1320 2358
rect 1280 2322 1284 2354
rect 1284 2322 1316 2354
rect 1316 2322 1320 2354
rect 1280 2318 1320 2322
rect 1192 2276 1232 2282
rect 1192 2244 1204 2276
rect 1204 2244 1232 2276
rect 1192 2242 1232 2244
rect -1588 1164 -1552 1184
rect 848 1722 888 1762
rect 1192 1758 1198 1772
rect 1198 1758 1230 1772
rect 1230 1758 1232 1772
rect 1192 1732 1232 1758
rect 936 1642 976 1660
rect 936 1620 940 1642
rect 940 1620 972 1642
rect 972 1620 976 1642
rect 1282 1716 1322 1720
rect 1282 1684 1286 1716
rect 1286 1684 1318 1716
rect 1318 1684 1322 1716
rect 1282 1680 1322 1684
rect -1074 720 -914 752
rect -1074 648 -914 720
rect -786 752 -626 758
rect -786 720 -626 752
rect -786 718 -626 720
rect -206 752 -46 756
rect -206 720 -46 752
rect -206 716 -46 720
rect 844 864 848 1242
rect 848 864 880 1242
rect 880 864 884 1242
rect 922 722 962 806
rect 1156 866 1160 1244
rect 1160 866 1192 1244
rect 1192 866 1196 1244
rect 1078 722 1118 806
rect 1000 300 1004 664
rect 1004 300 1036 664
rect 1036 300 1040 664
rect 1000 286 1040 300
rect 1234 722 1274 806
rect 1468 866 1472 1244
rect 1472 866 1504 1244
rect 1504 866 1508 1244
rect 1390 722 1430 806
rect 1312 300 1316 664
rect 1316 300 1348 664
rect 1348 300 1352 664
rect 1312 286 1352 300
rect 1546 722 1586 806
rect 1780 866 1784 1244
rect 1784 866 1816 1244
rect 1816 866 1820 1244
rect 1702 722 1742 806
rect 1624 300 1628 664
rect 1628 300 1660 664
rect 1660 300 1664 664
rect 1624 286 1664 300
rect 1858 722 1898 806
rect 2092 866 2096 1244
rect 2096 866 2128 1244
rect 2128 866 2132 1244
rect 2014 722 2054 806
rect 1936 300 1940 664
rect 1940 300 1972 664
rect 1972 300 1976 664
rect 1936 286 1976 300
rect 2170 722 2210 806
rect 2404 866 2408 1244
rect 2408 866 2440 1244
rect 2440 866 2444 1244
rect 2326 722 2366 806
rect 2248 300 2252 664
rect 2252 300 2284 664
rect 2284 300 2288 664
rect 2248 286 2288 300
rect -1682 -117 -1468 -94
rect -1682 -212 -1652 -117
rect -1652 -178 -1468 -117
rect -1652 -210 -1544 -178
rect -1544 -210 -1472 -178
rect -1472 -210 -1468 -178
rect -1652 -212 -1468 -210
rect 1656 -178 1888 -174
rect 1656 -210 1728 -178
rect 1728 -210 1816 -178
rect 1816 -210 1888 -178
rect 1656 -214 1888 -210
rect 2296 -178 2368 -174
rect 2296 -210 2368 -178
rect 2296 -214 2368 -210
rect -1680 -1182 -1652 -1090
rect -1652 -1122 -1544 -1090
rect -1544 -1122 -1472 -1090
rect -1472 -1122 -1466 -1090
rect -1652 -1182 -1466 -1122
rect -1680 -1208 -1466 -1182
<< metal2 >>
rect -1690 3026 -1458 3038
rect -1690 1164 -1592 3026
rect -1552 1164 -1458 3026
rect -1090 2832 38 2842
rect -1090 2498 -1080 2832
rect 28 2540 38 2832
rect 28 2498 742 2540
rect -1090 2488 742 2498
rect -16 2486 742 2488
rect 700 2410 742 2486
rect 700 2398 884 2410
rect 700 2358 836 2398
rect 876 2358 884 2398
rect 700 2344 884 2358
rect 1274 2358 1320 2368
rect 1274 2318 1280 2358
rect 914 2282 1232 2292
rect -300 2242 -8 2252
rect -300 2122 -290 2242
rect -1690 -94 -1458 1164
rect -1690 -212 -1682 -94
rect -1468 -212 -1458 -94
rect -1690 -1090 -1458 -212
rect -1362 2054 -742 2062
rect -1362 1944 -1074 2054
rect -760 1944 -742 2054
rect -1362 1934 -742 1944
rect -300 1938 -98 2122
rect -18 1938 -8 2242
rect 914 2242 924 2282
rect 964 2242 1192 2282
rect 914 2232 1232 2242
rect -1362 -182 -1196 1934
rect -300 1930 -8 1938
rect -256 1928 -8 1930
rect -250 1868 -78 1878
rect -1018 1828 -624 1868
rect -472 1828 -454 1868
rect -1018 1826 -454 1828
rect -250 1828 -240 1868
rect -88 1828 -78 1868
rect -1018 1770 -846 1826
rect -250 1776 -216 1828
rect -1018 1730 -1008 1770
rect -856 1730 -846 1770
rect -642 1774 -216 1776
rect -642 1734 -628 1774
rect -476 1734 -216 1774
rect -1018 766 -846 1730
rect -1092 752 -846 766
rect -250 1710 -216 1734
rect -114 1710 -78 1828
rect -250 1054 -78 1710
rect 544 1762 894 1782
rect 544 1722 848 1762
rect 888 1722 894 1762
rect 1192 1772 1232 2232
rect 1192 1722 1232 1732
rect 1274 1730 1320 2318
rect 544 1690 894 1722
rect 1274 1720 1328 1730
rect 544 1054 640 1690
rect 1274 1680 1282 1720
rect 1322 1680 1328 1720
rect 1274 1678 1328 1680
rect 936 1660 1328 1678
rect 976 1620 1328 1660
rect 936 1608 1328 1620
rect 736 1244 2554 1424
rect 736 1242 1156 1244
rect -250 944 642 1054
rect -250 762 -78 944
rect 532 806 642 944
rect 736 864 844 1242
rect 884 866 1156 1242
rect 1196 866 1468 1244
rect 1508 866 1780 1244
rect 1820 866 2092 1244
rect 2132 866 2404 1244
rect 2444 866 2554 1244
rect 884 864 2554 866
rect 736 854 2554 864
rect -1092 648 -1074 752
rect -914 648 -846 752
rect -800 758 -32 762
rect -800 718 -786 758
rect -626 756 -32 758
rect -626 718 -206 756
rect -800 716 -206 718
rect -46 716 -32 756
rect 532 722 922 806
rect 962 722 1078 806
rect 1118 722 1234 806
rect 1274 722 1390 806
rect 1430 722 1546 806
rect 1586 722 1702 806
rect 1742 722 1858 806
rect 1898 722 2014 806
rect 2054 722 2170 806
rect 2210 722 2326 806
rect 2366 722 2382 806
rect -800 668 -32 716
rect -1092 638 -846 648
rect 988 664 2562 674
rect 988 286 1000 664
rect 1040 286 1312 664
rect 1352 586 1624 664
rect 1664 586 1936 664
rect 1976 586 2248 664
rect 2288 586 2562 664
rect 1352 286 1528 586
rect 988 264 1528 286
rect 2326 264 2562 586
rect 988 74 2562 264
rect 1646 -174 1898 -164
rect 1646 -182 1656 -174
rect -1362 -214 1656 -182
rect 1888 -214 1898 -174
rect -1362 -224 1898 -214
rect 2282 -174 2382 74
rect 2282 -214 2296 -174
rect 2368 -214 2382 -174
rect 2282 -220 2382 -214
rect -1362 -328 1880 -224
rect -1690 -1208 -1680 -1090
rect -1466 -1208 -1458 -1090
rect -1690 -1218 -1458 -1208
<< via2 >>
rect -216 1710 -114 1828
rect 1528 286 1624 586
rect 1624 286 1664 586
rect 1664 286 1936 586
rect 1936 286 1976 586
rect 1976 286 2248 586
rect 2248 286 2288 586
rect 2288 286 2326 586
rect 1528 264 2326 286
<< metal3 >>
rect -626 1986 -300 1996
rect -626 1684 -616 1986
rect -256 1868 -246 1930
rect -256 1828 -86 1868
rect -256 1710 -216 1828
rect -114 1710 -86 1828
rect -256 1684 -86 1710
rect -626 1676 -86 1684
rect -626 1674 -246 1676
rect 1518 586 2336 596
rect 1518 264 1528 586
rect 2326 264 2336 586
rect 1518 254 2336 264
<< via3 >>
rect -616 1930 -300 1986
rect -616 1684 -256 1930
rect 1528 264 2326 586
<< metal4 >>
rect -626 1986 -246 1996
rect -626 1684 -616 1986
rect -256 1684 -246 1986
rect -626 1674 -246 1684
rect 1518 586 2336 596
rect 1518 264 1528 586
rect 2326 264 2336 586
rect 1518 254 2336 264
<< via4 >>
rect -616 1930 -300 1986
rect -300 1930 -256 1986
rect -616 1684 -256 1930
rect 1528 264 2326 586
<< metal5 >>
rect -694 1986 -168 2076
rect -694 1684 -616 1986
rect -256 1684 -168 1986
rect -694 1570 -168 1684
rect -1288 1450 952 1570
rect -1288 -550 -1168 1450
rect 832 -550 952 1450
rect 1518 586 2336 596
rect 1518 264 1528 586
rect 2326 264 2336 586
rect 1518 254 2336 264
rect -1288 -670 952 -550
<< via5 >>
rect 1528 264 2326 586
<< mimcapcontact >>
rect -1168 -550 832 1450
<< metal6 >>
rect -1288 1450 952 1570
rect -1288 -550 -1168 1450
rect 832 660 952 1450
rect 832 586 2414 660
rect 832 264 1528 586
rect 2326 264 2414 586
rect 832 182 2414 264
rect 832 -550 952 182
rect -1288 -670 952 -550
<< labels >>
flabel metal2 -1690 -94 -1458 1164 0 FreeSans 320 0 0 0 GND
port 2 nsew
flabel metal1 414 216 694 652 0 FreeSans 320 0 0 0 VCC
port 1 nsew
flabel metal2 -1090 2488 38 2842 1 FreeSans 320 0 0 0 ibias_1u
port 4 n
flabel metal2 1204 2036 1222 2098 1 FreeSans 320 0 0 0 en_n
port 6 n
flabel metal6 940 238 2362 638 0 FreeSans 320 0 0 0 out
port 5 nsew
flabel metal2 -288 1946 -48 2228 0 FreeSans 320 0 0 0 ref
port 3 nsew
<< end >>
