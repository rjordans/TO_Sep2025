magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754393324
<< nwell >>
rect -371 493 589 1463
rect -218 -843 149 -497
<< pwell >>
rect -286 -431 509 414
rect -267 -438 509 -431
rect 185 -529 509 -438
rect 195 -836 509 -529
rect 185 -837 509 -836
<< nmos >>
rect 221 -655 369 -629
<< pmos >>
rect -137 -655 87 -629
<< hvnmos >>
rect -90 211 310 301
rect -90 -139 310 -49
rect -90 -305 310 -215
<< hvpmos >>
rect -86 1099 -26 1189
rect 227 1099 287 1189
rect -90 841 310 921
rect -90 685 310 765
<< ndiff >>
rect 221 -575 369 -561
rect 221 -607 235 -575
rect 355 -607 369 -575
rect 221 -629 369 -607
rect 221 -677 369 -655
rect 221 -709 236 -677
rect 355 -709 369 -677
rect 221 -727 369 -709
<< pdiff >>
rect -137 -575 87 -559
rect -137 -607 -123 -575
rect 69 -607 87 -575
rect -137 -629 87 -607
rect -137 -677 87 -655
rect -137 -709 -119 -677
rect 70 -709 87 -677
rect -137 -731 87 -709
<< hvndiff >>
rect -90 355 310 369
rect -90 323 79 355
rect 296 323 310 355
rect -90 301 310 323
rect -90 189 310 211
rect -90 157 79 189
rect 296 157 310 189
rect -90 125 310 157
rect -90 5 310 23
rect -90 -27 -73 5
rect 25 -27 310 5
rect -90 -49 310 -27
rect -90 -161 310 -139
rect -90 -193 151 -161
rect 296 -193 310 -161
rect -90 -215 310 -193
rect -90 -327 310 -305
rect -90 -359 27 -327
rect 296 -359 310 -327
rect -90 -373 310 -359
<< hvpdiff >>
rect -86 1250 -26 1275
rect -86 1218 -72 1250
rect -40 1218 -26 1250
rect -86 1189 -26 1218
rect 227 1250 287 1275
rect 227 1218 241 1250
rect 273 1218 287 1250
rect 227 1189 287 1218
rect -86 1077 -26 1099
rect -86 1045 -72 1077
rect -40 1045 -26 1077
rect -86 1031 -26 1045
rect 227 1077 287 1099
rect 227 1045 241 1077
rect 273 1045 287 1077
rect 227 1031 287 1045
rect -90 975 310 989
rect -90 943 9 975
rect 296 943 310 975
rect -90 921 310 943
rect -90 819 310 841
rect -90 787 120 819
rect 296 787 310 819
rect -90 765 310 787
rect -90 663 310 685
rect -90 631 6 663
rect 296 631 310 663
rect -90 617 310 631
<< ndiffc >>
rect 235 -607 355 -575
rect 236 -709 355 -677
<< pdiffc >>
rect -123 -607 69 -575
rect -119 -709 70 -677
<< hvndiffc >>
rect 79 323 296 355
rect 79 157 296 189
rect -73 -27 25 5
rect 151 -193 296 -161
rect 27 -359 296 -327
<< hvpdiffc >>
rect -72 1218 -40 1250
rect 241 1218 273 1250
rect -72 1045 -40 1077
rect 241 1045 273 1077
rect 9 943 296 975
rect 120 787 296 819
rect 6 631 296 663
<< psubdiff >>
rect 221 -745 369 -727
rect 221 -777 236 -745
rect 355 -777 369 -745
rect 221 -791 369 -777
<< nsubdiff >>
rect -137 -749 87 -731
rect -137 -781 -119 -749
rect 70 -781 87 -749
rect -137 -795 87 -781
<< hvpsubdiff >>
rect -246 355 -186 369
rect -246 -359 -232 355
rect -200 125 -186 355
rect 405 355 465 369
rect 405 125 419 355
rect -200 65 419 125
rect -200 -359 -186 65
rect -246 -373 -186 -359
rect 405 -365 419 65
rect 451 -365 465 355
rect 405 -379 465 -365
<< hvnsubdiff >>
rect -246 1325 465 1339
rect -246 631 -232 1325
rect -200 1293 -164 1325
rect -108 1293 -4 1325
rect 205 1293 309 1325
rect 383 1293 419 1325
rect -200 1275 419 1293
rect -200 631 -186 1275
rect -246 617 -186 631
rect 405 631 419 1275
rect 451 631 465 1325
rect 405 617 465 631
<< psubdiffcont >>
rect 236 -777 355 -745
<< nsubdiffcont >>
rect -119 -781 70 -749
<< hvpsubdiffcont >>
rect -232 -359 -200 355
rect 419 -365 451 355
<< hvnsubdiffcont >>
rect -232 631 -200 1325
rect -164 1293 -108 1325
rect -4 1293 205 1325
rect 309 1293 383 1325
rect 419 631 451 1325
<< poly >>
rect -164 1167 -86 1189
rect -164 1116 -150 1167
rect -118 1116 -86 1167
rect -164 1099 -86 1116
rect -26 1099 10 1189
rect 105 1099 227 1189
rect 287 1099 323 1189
rect 105 1089 207 1099
rect 105 1017 120 1089
rect 193 1017 207 1089
rect 105 1003 207 1017
rect -164 907 -90 921
rect -164 856 -150 907
rect -118 856 -90 907
rect -164 841 -90 856
rect 310 841 355 921
rect -164 765 -112 841
rect -164 751 -90 765
rect -164 700 -150 751
rect -118 700 -90 751
rect -164 685 -90 700
rect 310 685 355 765
rect -164 301 -112 685
rect -164 287 -90 301
rect -164 225 -150 287
rect -118 225 -90 287
rect -164 211 -90 225
rect 310 211 346 301
rect -164 -63 -90 -49
rect -164 -125 -150 -63
rect -118 -125 -90 -63
rect -164 -139 -90 -125
rect 310 -139 346 -49
rect -164 -229 -90 -215
rect -164 -291 -150 -229
rect -118 -291 -90 -229
rect -164 -305 -90 -291
rect 310 -305 346 -215
rect 110 -469 170 -455
rect 110 -501 124 -469
rect 156 -501 170 -469
rect 110 -515 170 -501
rect 127 -629 153 -515
rect -173 -655 -137 -629
rect 87 -655 221 -629
rect 369 -655 405 -629
<< polycont >>
rect -150 1116 -118 1167
rect 120 1017 193 1089
rect -150 856 -118 907
rect -150 700 -118 751
rect -150 225 -118 287
rect -150 -125 -118 -63
rect -150 -291 -118 -229
rect 124 -501 156 -469
<< metal1 >>
rect -246 1325 465 1339
rect -246 631 -232 1325
rect -200 1293 -164 1325
rect -108 1293 -4 1325
rect 205 1293 309 1325
rect 383 1293 419 1325
rect -200 1250 419 1293
rect -200 1219 -72 1250
rect -200 631 -186 1219
rect -82 1218 -72 1219
rect -40 1218 241 1250
rect 273 1218 419 1250
rect -246 617 -186 631
rect -150 1167 -118 1177
rect -118 1125 273 1158
rect -150 907 -118 1116
rect -150 751 -118 856
rect -246 355 -186 369
rect -246 -359 -232 355
rect -200 -359 -186 355
rect -150 287 -118 700
rect -73 1077 -38 1089
rect 106 1077 120 1089
rect -73 1045 -72 1077
rect -40 1045 120 1077
rect -73 353 -38 1045
rect 106 1017 120 1045
rect 193 1017 205 1089
rect 241 1077 273 1125
rect 241 1034 273 1045
rect -2 943 9 975
rect 296 943 311 975
rect 6 673 73 943
rect 405 819 419 1218
rect 109 787 120 819
rect 296 787 419 819
rect 6 663 296 673
rect 6 400 296 631
rect 405 631 419 787
rect 451 631 465 1325
rect 405 616 465 631
rect 79 355 296 400
rect -73 318 33 353
rect -118 235 -40 267
rect -150 214 -118 225
rect -73 16 -40 235
rect -2 98 33 318
rect 79 313 296 323
rect 405 355 465 369
rect 405 189 419 355
rect 69 157 79 189
rect 296 157 419 189
rect -2 63 105 98
rect -73 5 25 16
rect -73 -37 25 -27
rect -150 -63 -118 -53
rect -118 -115 -9 -83
rect -150 -136 -118 -125
rect -246 -373 -186 -359
rect -150 -229 -118 -215
rect -150 -564 -118 -291
rect -41 -469 -9 -115
rect 70 -312 105 63
rect 405 -161 419 157
rect 141 -193 151 -161
rect 296 -193 419 -161
rect 27 -327 296 -312
rect 27 -377 296 -359
rect 405 -365 419 -193
rect 451 -365 465 355
rect -41 -501 124 -469
rect 156 -501 166 -469
rect -150 -575 369 -564
rect -150 -607 -123 -575
rect 69 -607 235 -575
rect 355 -607 369 -575
rect -150 -617 369 -607
rect 405 -667 465 -365
rect -119 -677 70 -667
rect -119 -749 70 -709
rect -119 -791 70 -781
rect 236 -677 465 -667
rect 355 -709 465 -677
rect 236 -745 465 -709
rect 355 -777 465 -745
rect 236 -787 465 -777
<< labels >>
flabel hvpsubdiffcont 429 -182 434 -167 1 FreeSans 320 0 0 0 GND
port 3 n power default
flabel metal1 -133 -346 -133 -346 1 FreeSans 320 0 0 0 in_b
flabel hvpsubdiffcont -222 -182 -217 -167 1 FreeSans 320 0 0 0 GND
flabel metal1 -29 -723 -29 -723 0 FreeSans 320 0 0 0 VDD_1v2
port 2 nsew power default
flabel metal1 58 -490 58 -490 0 FreeSans 320 0 0 0 in
port 4 nsew
flabel hvndiffc 110 -349 110 -349 0 FreeSans 320 0 0 0 lvlsh
flabel hvndiffc -26 -16 -26 -16 0 FreeSans 320 0 0 0 lvlsh_b
flabel metal1 183 482 183 482 1 FreeSans 320 0 0 0 out
port 5 n
flabel hvnsubdiffcont 74 1319 74 1319 0 FreeSans 320 0 0 0 VDD_3v3
port 1 nsew power default
<< end >>
