magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757254581
<< nwell >>
rect 5172 3297 6176 5505
rect 3170 1948 6112 2580
rect 4038 1146 6112 1948
rect 3132 6 6112 1146
<< hvnmos >>
rect 3300 5063 3700 5263
rect 3878 5063 4278 5263
rect 4456 5063 4856 5263
rect 3300 4679 3700 4879
rect 3878 4679 4278 4879
rect 4456 4679 4856 4879
rect 3300 4295 3700 4495
rect 3878 4295 4278 4495
rect 4456 4295 4856 4495
rect 3300 3911 3700 4111
rect 3878 3911 4278 4111
rect 4456 3911 4856 4111
rect 3300 3527 3700 3727
rect 3878 3527 4278 3727
rect 4456 3527 4856 3727
rect 3458 2872 3548 2932
rect 3734 2872 3824 2932
<< hvpmos >>
rect 5470 5027 5870 5227
rect 5470 4739 5870 4939
rect 5470 4451 5870 4651
rect 5470 4163 5870 4363
rect 5470 3875 5870 4075
rect 5470 3587 5870 3787
rect 3476 2234 3556 2294
rect 3734 2234 3814 2294
rect 3402 770 3802 850
rect 3402 614 3802 694
rect 3402 458 3802 538
rect 3402 302 3802 382
rect 4332 292 4412 2292
rect 4488 292 4568 2292
rect 4644 292 4724 2292
rect 4800 292 4880 2292
rect 4956 292 5036 2292
rect 5112 292 5192 2292
rect 5268 292 5348 2292
rect 5424 292 5504 2292
rect 5580 292 5660 2292
rect 5736 292 5816 2292
<< hvndiff >>
rect 3232 5249 3300 5263
rect 3232 5077 3246 5249
rect 3278 5077 3300 5249
rect 3232 5063 3300 5077
rect 3700 5249 3768 5263
rect 3700 5077 3722 5249
rect 3754 5077 3768 5249
rect 3700 5063 3768 5077
rect 3810 5249 3878 5263
rect 3810 5077 3824 5249
rect 3856 5077 3878 5249
rect 3810 5063 3878 5077
rect 4278 5249 4346 5263
rect 4278 5077 4300 5249
rect 4332 5077 4346 5249
rect 4278 5063 4346 5077
rect 4388 5249 4456 5263
rect 4388 5077 4402 5249
rect 4434 5077 4456 5249
rect 4388 5063 4456 5077
rect 4856 5249 4924 5263
rect 4856 5077 4878 5249
rect 4910 5077 4924 5249
rect 4856 5063 4924 5077
rect 3232 4865 3300 4879
rect 3232 4693 3246 4865
rect 3278 4693 3300 4865
rect 3232 4679 3300 4693
rect 3700 4865 3768 4879
rect 3700 4693 3722 4865
rect 3754 4693 3768 4865
rect 3700 4679 3768 4693
rect 3810 4865 3878 4879
rect 3810 4693 3824 4865
rect 3856 4693 3878 4865
rect 3810 4679 3878 4693
rect 4278 4865 4346 4879
rect 4278 4693 4300 4865
rect 4332 4693 4346 4865
rect 4278 4679 4346 4693
rect 4388 4865 4456 4879
rect 4388 4693 4402 4865
rect 4434 4693 4456 4865
rect 4388 4679 4456 4693
rect 4856 4865 4924 4879
rect 4856 4693 4878 4865
rect 4910 4693 4924 4865
rect 4856 4679 4924 4693
rect 3232 4481 3300 4495
rect 3232 4309 3246 4481
rect 3278 4309 3300 4481
rect 3232 4295 3300 4309
rect 3700 4481 3768 4495
rect 3700 4309 3722 4481
rect 3754 4309 3768 4481
rect 3700 4295 3768 4309
rect 3810 4481 3878 4495
rect 3810 4309 3824 4481
rect 3856 4309 3878 4481
rect 3810 4295 3878 4309
rect 4278 4481 4346 4495
rect 4278 4309 4300 4481
rect 4332 4309 4346 4481
rect 4278 4295 4346 4309
rect 4388 4481 4456 4495
rect 4388 4309 4402 4481
rect 4434 4309 4456 4481
rect 4388 4295 4456 4309
rect 4856 4481 4924 4495
rect 4856 4309 4878 4481
rect 4910 4309 4924 4481
rect 4856 4295 4924 4309
rect 3232 4097 3300 4111
rect 3232 3925 3246 4097
rect 3278 3925 3300 4097
rect 3232 3911 3300 3925
rect 3700 4097 3768 4111
rect 3700 3925 3722 4097
rect 3754 3925 3768 4097
rect 3700 3911 3768 3925
rect 3810 4097 3878 4111
rect 3810 3925 3824 4097
rect 3856 3925 3878 4097
rect 3810 3911 3878 3925
rect 4278 4097 4346 4111
rect 4278 3925 4300 4097
rect 4332 3925 4346 4097
rect 4278 3911 4346 3925
rect 4388 4097 4456 4111
rect 4388 3925 4402 4097
rect 4434 3925 4456 4097
rect 4388 3911 4456 3925
rect 4856 4097 4924 4111
rect 4856 3925 4878 4097
rect 4910 3925 4924 4097
rect 4856 3911 4924 3925
rect 3232 3713 3300 3727
rect 3232 3541 3246 3713
rect 3278 3541 3300 3713
rect 3232 3527 3300 3541
rect 3700 3713 3768 3727
rect 3700 3541 3722 3713
rect 3754 3541 3768 3713
rect 3700 3527 3768 3541
rect 3810 3713 3878 3727
rect 3810 3541 3824 3713
rect 3856 3541 3878 3713
rect 3810 3527 3878 3541
rect 4278 3713 4346 3727
rect 4278 3541 4300 3713
rect 4332 3541 4346 3713
rect 4278 3527 4346 3541
rect 4388 3713 4456 3727
rect 4388 3541 4402 3713
rect 4434 3541 4456 3713
rect 4388 3527 4456 3541
rect 4856 3713 4924 3727
rect 4856 3541 4878 3713
rect 4910 3541 4924 3713
rect 4856 3527 4924 3541
rect 3390 2918 3458 2932
rect 3390 2886 3404 2918
rect 3436 2886 3458 2918
rect 3390 2872 3458 2886
rect 3548 2918 3734 2932
rect 3548 2886 3570 2918
rect 3712 2886 3734 2918
rect 3548 2872 3734 2886
rect 3824 2918 3892 2932
rect 3824 2886 3846 2918
rect 3878 2886 3892 2918
rect 3824 2872 3892 2886
<< hvpdiff >>
rect 5398 5213 5470 5227
rect 5398 5041 5416 5213
rect 5448 5041 5470 5213
rect 5398 5027 5470 5041
rect 5870 5213 5948 5227
rect 5870 5041 5902 5213
rect 5934 5041 5948 5213
rect 5870 5027 5948 5041
rect 5398 4925 5470 4939
rect 5398 4753 5416 4925
rect 5448 4753 5470 4925
rect 5398 4739 5470 4753
rect 5870 4925 5948 4939
rect 5870 4753 5902 4925
rect 5934 4753 5948 4925
rect 5870 4739 5948 4753
rect 5398 4637 5470 4651
rect 5398 4465 5416 4637
rect 5448 4465 5470 4637
rect 5398 4451 5470 4465
rect 5870 4637 5948 4651
rect 5870 4465 5902 4637
rect 5934 4465 5948 4637
rect 5870 4451 5948 4465
rect 5398 4349 5470 4363
rect 5398 4177 5416 4349
rect 5448 4177 5470 4349
rect 5398 4163 5470 4177
rect 5870 4349 5948 4363
rect 5870 4177 5902 4349
rect 5934 4177 5948 4349
rect 5870 4163 5948 4177
rect 5398 4061 5470 4075
rect 5398 3889 5416 4061
rect 5448 3889 5470 4061
rect 5398 3875 5470 3889
rect 5870 4061 5948 4075
rect 5870 3889 5902 4061
rect 5934 3889 5948 4061
rect 5870 3875 5948 3889
rect 5398 3773 5470 3787
rect 5398 3601 5416 3773
rect 5448 3601 5470 3773
rect 5398 3587 5470 3601
rect 5870 3773 5946 3787
rect 5870 3601 5900 3773
rect 5932 3601 5946 3773
rect 5870 3587 5946 3601
rect 3408 2280 3476 2294
rect 3408 2248 3422 2280
rect 3454 2248 3476 2280
rect 3408 2234 3476 2248
rect 3556 2280 3734 2294
rect 3556 2248 3582 2280
rect 3712 2248 3734 2280
rect 3556 2234 3734 2248
rect 3814 2280 3894 2294
rect 3814 2248 3848 2280
rect 3880 2248 3894 2280
rect 3814 2234 3894 2248
rect 3402 904 3802 918
rect 3402 872 3416 904
rect 3788 872 3802 904
rect 3402 850 3802 872
rect 3402 748 3802 770
rect 3402 716 3416 748
rect 3788 716 3802 748
rect 3402 694 3802 716
rect 3402 592 3802 614
rect 3402 560 3416 592
rect 3788 560 3802 592
rect 3402 538 3802 560
rect 3402 436 3802 458
rect 3402 404 3416 436
rect 3788 404 3802 436
rect 3402 382 3802 404
rect 3402 280 3802 302
rect 3402 248 3416 280
rect 3788 248 3802 280
rect 3402 234 3802 248
rect 4264 2268 4332 2292
rect 4264 312 4278 2268
rect 4310 312 4332 2268
rect 4264 292 4332 312
rect 4412 2270 4488 2292
rect 4412 314 4434 2270
rect 4466 314 4488 2270
rect 4412 292 4488 314
rect 4568 2270 4644 2292
rect 4568 314 4590 2270
rect 4622 314 4644 2270
rect 4568 292 4644 314
rect 4724 2270 4800 2292
rect 4724 314 4746 2270
rect 4778 314 4800 2270
rect 4724 292 4800 314
rect 4880 2270 4956 2292
rect 4880 314 4902 2270
rect 4934 314 4956 2270
rect 4880 292 4956 314
rect 5036 2270 5112 2292
rect 5036 314 5058 2270
rect 5090 314 5112 2270
rect 5036 292 5112 314
rect 5192 2270 5268 2292
rect 5192 314 5214 2270
rect 5246 314 5268 2270
rect 5192 292 5268 314
rect 5348 2270 5424 2292
rect 5348 314 5370 2270
rect 5402 314 5424 2270
rect 5348 292 5424 314
rect 5504 2270 5580 2292
rect 5504 314 5526 2270
rect 5558 314 5580 2270
rect 5504 292 5580 314
rect 5660 2270 5736 2292
rect 5660 314 5682 2270
rect 5714 314 5736 2270
rect 5660 292 5736 314
rect 5816 2270 5884 2292
rect 5816 314 5838 2270
rect 5870 314 5884 2270
rect 5816 292 5884 314
<< hvndiffc >>
rect 3246 5077 3278 5249
rect 3722 5077 3754 5249
rect 3824 5077 3856 5249
rect 4300 5077 4332 5249
rect 4402 5077 4434 5249
rect 4878 5077 4910 5249
rect 3246 4693 3278 4865
rect 3722 4693 3754 4865
rect 3824 4693 3856 4865
rect 4300 4693 4332 4865
rect 4402 4693 4434 4865
rect 4878 4693 4910 4865
rect 3246 4309 3278 4481
rect 3722 4309 3754 4481
rect 3824 4309 3856 4481
rect 4300 4309 4332 4481
rect 4402 4309 4434 4481
rect 4878 4309 4910 4481
rect 3246 3925 3278 4097
rect 3722 3925 3754 4097
rect 3824 3925 3856 4097
rect 4300 3925 4332 4097
rect 4402 3925 4434 4097
rect 4878 3925 4910 4097
rect 3246 3541 3278 3713
rect 3722 3541 3754 3713
rect 3824 3541 3856 3713
rect 4300 3541 4332 3713
rect 4402 3541 4434 3713
rect 4878 3541 4910 3713
rect 3404 2886 3436 2918
rect 3570 2886 3712 2918
rect 3846 2886 3878 2918
<< hvpdiffc >>
rect 5416 5041 5448 5213
rect 5902 5041 5934 5213
rect 5416 4753 5448 4925
rect 5902 4753 5934 4925
rect 5416 4465 5448 4637
rect 5902 4465 5934 4637
rect 5416 4177 5448 4349
rect 5902 4177 5934 4349
rect 5416 3889 5448 4061
rect 5902 3889 5934 4061
rect 5416 3601 5448 3773
rect 5900 3601 5932 3773
rect 3422 2248 3454 2280
rect 3582 2248 3712 2280
rect 3848 2248 3880 2280
rect 3416 872 3788 904
rect 3416 716 3788 748
rect 3416 560 3788 592
rect 3416 404 3788 436
rect 3416 248 3788 280
rect 4278 312 4310 2268
rect 4434 314 4466 2270
rect 4590 314 4622 2270
rect 4746 314 4778 2270
rect 4902 314 4934 2270
rect 5058 314 5090 2270
rect 5214 314 5246 2270
rect 5370 314 5402 2270
rect 5526 314 5558 2270
rect 5682 314 5714 2270
rect 5838 314 5870 2270
<< psubdiff >>
rect -14 5435 3084 5449
rect -14 10 0 5435
rect 32 5389 3038 5403
rect 32 56 46 5389
rect 3024 56 3038 5389
rect 32 42 3038 56
rect 3070 10 3084 5435
rect -14 -4 3084 10
<< hvpsubdiff >>
rect 3128 5435 5030 5449
rect 3128 3381 3142 5435
rect 3174 5389 4984 5403
rect 3174 3427 3188 5389
rect 4970 3427 4984 5389
rect 3174 3413 4984 3427
rect 5016 3381 5030 5435
rect 3128 3367 5030 3381
rect 3288 3090 3994 3104
rect 3288 2718 3302 3090
rect 3334 3044 3948 3058
rect 3334 2764 3348 3044
rect 3934 2764 3948 3044
rect 3334 2750 3948 2764
rect 3980 2718 3994 3090
rect 3288 2704 3994 2718
<< hvnsubdiff >>
rect 5296 5367 6052 5381
rect 5296 3435 5310 5367
rect 5342 5313 6006 5335
rect 5342 3489 5356 5313
rect 5992 3489 6006 5313
rect 5342 3467 6006 3489
rect 6038 3435 6052 5367
rect 5296 3421 6052 3435
rect 3306 2442 3996 2456
rect 3306 2086 3320 2442
rect 3352 2396 3950 2410
rect 3352 2132 3366 2396
rect 3936 2132 3950 2396
rect 3352 2118 3950 2132
rect 3982 2086 3996 2442
rect 3306 2072 3996 2086
rect 4162 2442 5988 2456
rect 3256 1006 4036 1020
rect 3256 146 3270 1006
rect 3302 960 3990 974
rect 3302 192 3316 960
rect 3976 192 3990 960
rect 3302 178 3990 192
rect 4022 146 4036 1006
rect 3256 132 4036 146
rect 4162 144 4176 2442
rect 4208 2396 5942 2410
rect 4208 190 4222 2396
rect 5928 190 5942 2396
rect 4208 176 5942 190
rect 5974 144 5988 2442
rect 4162 130 5988 144
<< psubdiffcont >>
rect 0 5403 3070 5435
rect 0 42 32 5403
rect 3038 42 3070 5403
rect 0 10 3070 42
<< hvpsubdiffcont >>
rect 3142 5403 5016 5435
rect 3142 3413 3174 5403
rect 4984 3413 5016 5403
rect 3142 3381 5016 3413
rect 3302 3058 3980 3090
rect 3302 2750 3334 3058
rect 3948 2750 3980 3058
rect 3302 2718 3980 2750
<< hvnsubdiffcont >>
rect 5310 5335 6038 5367
rect 5310 3467 5342 5335
rect 6006 3467 6038 5335
rect 5310 3435 6038 3467
rect 3320 2410 3982 2442
rect 3320 2118 3352 2410
rect 3950 2118 3982 2410
rect 3320 2086 3982 2118
rect 3270 974 4022 1006
rect 3270 178 3302 974
rect 3990 178 4022 974
rect 3270 146 4022 178
rect 4176 2410 5974 2442
rect 4176 176 4208 2410
rect 5942 176 5974 2410
rect 4176 144 5974 176
<< poly >>
rect 126 5343 226 5357
rect 126 5311 140 5343
rect 212 5311 226 5343
rect 126 5271 226 5311
rect 126 2831 226 2871
rect 126 2799 140 2831
rect 212 2799 226 2831
rect 126 2785 226 2799
rect 286 5343 386 5357
rect 286 5311 300 5343
rect 372 5311 386 5343
rect 286 5271 386 5311
rect 286 2831 386 2871
rect 286 2799 300 2831
rect 372 2799 386 2831
rect 286 2785 386 2799
rect 446 5343 546 5357
rect 446 5311 460 5343
rect 532 5311 546 5343
rect 446 5271 546 5311
rect 446 2831 546 2871
rect 446 2799 460 2831
rect 532 2799 546 2831
rect 446 2785 546 2799
rect 606 5343 706 5357
rect 606 5311 620 5343
rect 692 5311 706 5343
rect 606 5271 706 5311
rect 606 2831 706 2871
rect 606 2799 620 2831
rect 692 2799 706 2831
rect 606 2785 706 2799
rect 766 5343 866 5357
rect 766 5311 780 5343
rect 852 5311 866 5343
rect 766 5271 866 5311
rect 766 2831 866 2871
rect 766 2799 780 2831
rect 852 2799 866 2831
rect 766 2785 866 2799
rect 926 5343 1026 5357
rect 926 5311 940 5343
rect 1012 5311 1026 5343
rect 926 5271 1026 5311
rect 926 2831 1026 2871
rect 926 2799 940 2831
rect 1012 2799 1026 2831
rect 926 2785 1026 2799
rect 1086 5343 1186 5357
rect 1086 5311 1100 5343
rect 1172 5311 1186 5343
rect 1086 5271 1186 5311
rect 1086 2831 1186 2871
rect 1086 2799 1100 2831
rect 1172 2799 1186 2831
rect 1086 2785 1186 2799
rect 1246 5343 1346 5357
rect 1246 5311 1260 5343
rect 1332 5311 1346 5343
rect 1246 5271 1346 5311
rect 1246 2831 1346 2871
rect 1246 2799 1260 2831
rect 1332 2799 1346 2831
rect 1246 2785 1346 2799
rect 1406 5343 1506 5357
rect 1406 5311 1420 5343
rect 1492 5311 1506 5343
rect 1406 5271 1506 5311
rect 1406 2831 1506 2871
rect 1406 2799 1420 2831
rect 1492 2799 1506 2831
rect 1406 2785 1506 2799
rect 1566 5343 1666 5357
rect 1566 5311 1580 5343
rect 1652 5311 1666 5343
rect 1566 5271 1666 5311
rect 1566 2831 1666 2871
rect 1566 2799 1580 2831
rect 1652 2799 1666 2831
rect 1566 2785 1666 2799
rect 1726 5343 1826 5357
rect 1726 5311 1740 5343
rect 1812 5311 1826 5343
rect 1726 5271 1826 5311
rect 1726 2831 1826 2871
rect 1726 2799 1740 2831
rect 1812 2799 1826 2831
rect 1726 2785 1826 2799
rect 1886 5343 1986 5357
rect 1886 5311 1900 5343
rect 1972 5311 1986 5343
rect 1886 5271 1986 5311
rect 1886 2831 1986 2871
rect 1886 2799 1900 2831
rect 1972 2799 1986 2831
rect 1886 2785 1986 2799
rect 2046 5343 2146 5357
rect 2046 5311 2060 5343
rect 2132 5311 2146 5343
rect 2046 5271 2146 5311
rect 2046 2831 2146 2871
rect 2046 2799 2060 2831
rect 2132 2799 2146 2831
rect 2046 2785 2146 2799
rect 2206 5343 2306 5357
rect 2206 5311 2220 5343
rect 2292 5311 2306 5343
rect 2206 5271 2306 5311
rect 2206 2831 2306 2871
rect 2206 2799 2220 2831
rect 2292 2799 2306 2831
rect 2206 2785 2306 2799
rect 2366 5343 2466 5357
rect 2366 5311 2380 5343
rect 2452 5311 2466 5343
rect 2366 5271 2466 5311
rect 2366 2831 2466 2871
rect 2366 2799 2380 2831
rect 2452 2799 2466 2831
rect 2366 2785 2466 2799
rect 2526 5343 2626 5357
rect 2526 5311 2540 5343
rect 2612 5311 2626 5343
rect 2526 5271 2626 5311
rect 2526 2831 2626 2871
rect 2526 2799 2540 2831
rect 2612 2799 2626 2831
rect 2526 2785 2626 2799
rect 2686 5343 2786 5357
rect 2686 5311 2700 5343
rect 2772 5311 2786 5343
rect 2686 5271 2786 5311
rect 2686 2831 2786 2871
rect 2686 2799 2700 2831
rect 2772 2799 2786 2831
rect 2686 2785 2786 2799
rect 2844 5343 2944 5357
rect 2844 5311 2858 5343
rect 2930 5311 2944 5343
rect 2844 5271 2944 5311
rect 2844 2831 2944 2871
rect 2844 2799 2858 2831
rect 2930 2799 2944 2831
rect 2844 2785 2944 2799
rect 126 2647 226 2661
rect 126 2615 140 2647
rect 212 2615 226 2647
rect 126 2575 226 2615
rect 126 135 226 175
rect 126 103 140 135
rect 212 103 226 135
rect 126 89 226 103
rect 286 2647 386 2661
rect 286 2615 300 2647
rect 372 2615 386 2647
rect 286 2575 386 2615
rect 286 135 386 175
rect 286 103 300 135
rect 372 103 386 135
rect 286 89 386 103
rect 446 2647 546 2661
rect 446 2615 460 2647
rect 532 2615 546 2647
rect 446 2575 546 2615
rect 446 135 546 175
rect 446 103 460 135
rect 532 103 546 135
rect 446 89 546 103
rect 606 2647 706 2661
rect 606 2615 620 2647
rect 692 2615 706 2647
rect 606 2575 706 2615
rect 606 135 706 175
rect 606 103 620 135
rect 692 103 706 135
rect 606 89 706 103
rect 766 2647 866 2661
rect 766 2615 780 2647
rect 852 2615 866 2647
rect 766 2575 866 2615
rect 766 135 866 175
rect 766 103 780 135
rect 852 103 866 135
rect 766 89 866 103
rect 926 2647 1026 2661
rect 926 2615 940 2647
rect 1012 2615 1026 2647
rect 926 2575 1026 2615
rect 926 135 1026 175
rect 926 103 940 135
rect 1012 103 1026 135
rect 926 89 1026 103
rect 1086 2647 1186 2661
rect 1086 2615 1100 2647
rect 1172 2615 1186 2647
rect 1086 2575 1186 2615
rect 1086 135 1186 175
rect 1086 103 1100 135
rect 1172 103 1186 135
rect 1086 89 1186 103
rect 1246 2647 1346 2661
rect 1246 2615 1260 2647
rect 1332 2615 1346 2647
rect 1246 2575 1346 2615
rect 1246 135 1346 175
rect 1246 103 1260 135
rect 1332 103 1346 135
rect 1246 89 1346 103
rect 1406 2647 1506 2661
rect 1406 2615 1420 2647
rect 1492 2615 1506 2647
rect 1406 2575 1506 2615
rect 1406 135 1506 175
rect 1406 103 1420 135
rect 1492 103 1506 135
rect 1406 89 1506 103
rect 1566 2647 1666 2661
rect 1566 2615 1580 2647
rect 1652 2615 1666 2647
rect 1566 2575 1666 2615
rect 1566 135 1666 175
rect 1566 103 1580 135
rect 1652 103 1666 135
rect 1566 89 1666 103
rect 1726 2647 1826 2661
rect 1726 2615 1740 2647
rect 1812 2615 1826 2647
rect 1726 2575 1826 2615
rect 1726 135 1826 175
rect 1726 103 1740 135
rect 1812 103 1826 135
rect 1726 89 1826 103
rect 1886 2647 1986 2661
rect 1886 2615 1900 2647
rect 1972 2615 1986 2647
rect 1886 2575 1986 2615
rect 1886 135 1986 175
rect 1886 103 1900 135
rect 1972 103 1986 135
rect 1886 89 1986 103
rect 2046 2647 2146 2661
rect 2046 2615 2060 2647
rect 2132 2615 2146 2647
rect 2046 2575 2146 2615
rect 2046 135 2146 175
rect 2046 103 2060 135
rect 2132 103 2146 135
rect 2046 89 2146 103
rect 2206 2647 2306 2661
rect 2206 2615 2220 2647
rect 2292 2615 2306 2647
rect 2206 2575 2306 2615
rect 2206 135 2306 175
rect 2206 103 2220 135
rect 2292 103 2306 135
rect 2206 89 2306 103
rect 2366 2647 2466 2661
rect 2366 2615 2380 2647
rect 2452 2615 2466 2647
rect 2366 2575 2466 2615
rect 2366 135 2466 175
rect 2366 103 2380 135
rect 2452 103 2466 135
rect 2366 89 2466 103
rect 2526 2647 2626 2661
rect 2526 2615 2540 2647
rect 2612 2615 2626 2647
rect 2526 2575 2626 2615
rect 2526 135 2626 175
rect 2526 103 2540 135
rect 2612 103 2626 135
rect 2526 89 2626 103
rect 2686 2647 2786 2661
rect 2686 2615 2700 2647
rect 2772 2615 2786 2647
rect 2686 2575 2786 2615
rect 2686 135 2786 175
rect 2686 103 2700 135
rect 2772 103 2786 135
rect 2686 89 2786 103
rect 2844 2647 2944 2661
rect 2844 2615 2858 2647
rect 2930 2615 2944 2647
rect 2844 2575 2944 2615
rect 2844 135 2944 175
rect 2844 103 2858 135
rect 2930 103 2944 135
rect 2844 89 2944 103
rect 3300 5323 3700 5337
rect 3300 5291 3324 5323
rect 3686 5291 3700 5323
rect 3300 5263 3700 5291
rect 3878 5323 4278 5337
rect 3878 5291 3902 5323
rect 4264 5291 4278 5323
rect 3878 5263 4278 5291
rect 4456 5323 4856 5337
rect 4456 5291 4470 5323
rect 4832 5291 4856 5323
rect 4456 5263 4856 5291
rect 3300 5035 3700 5063
rect 3300 5003 3324 5035
rect 3686 5003 3700 5035
rect 3300 4989 3700 5003
rect 3878 5035 4278 5063
rect 3878 5003 3902 5035
rect 4264 5003 4278 5035
rect 3878 4989 4278 5003
rect 4456 5035 4856 5063
rect 4456 5003 4470 5035
rect 4832 5003 4856 5035
rect 4456 4989 4856 5003
rect 3300 4939 3700 4953
rect 3300 4907 3334 4939
rect 3666 4907 3700 4939
rect 3300 4879 3700 4907
rect 3878 4939 4278 4953
rect 3878 4907 3902 4939
rect 4056 4907 4278 4939
rect 3878 4879 4278 4907
rect 4456 4939 4856 4953
rect 4456 4907 4470 4939
rect 4832 4907 4856 4939
rect 4456 4879 4856 4907
rect 3300 4651 3700 4679
rect 3300 4619 3334 4651
rect 3666 4619 3700 4651
rect 3300 4605 3700 4619
rect 3878 4651 4278 4679
rect 3878 4619 3902 4651
rect 4056 4619 4278 4651
rect 3878 4605 4278 4619
rect 4456 4651 4856 4679
rect 4456 4619 4490 4651
rect 4832 4619 4856 4651
rect 4456 4605 4856 4619
rect 3300 4555 3700 4569
rect 3300 4523 3334 4555
rect 3666 4523 3700 4555
rect 3300 4495 3700 4523
rect 3878 4555 4278 4569
rect 3878 4523 4100 4555
rect 4254 4523 4278 4555
rect 3878 4495 4278 4523
rect 4456 4555 4856 4569
rect 4456 4523 4480 4555
rect 4634 4523 4856 4555
rect 4456 4495 4856 4523
rect 3300 4267 3700 4295
rect 3300 4235 3334 4267
rect 3666 4235 3700 4267
rect 3300 4221 3700 4235
rect 3878 4267 4278 4295
rect 3878 4235 4100 4267
rect 4254 4235 4278 4267
rect 3878 4221 4278 4235
rect 4456 4267 4856 4295
rect 4456 4235 4480 4267
rect 4634 4235 4856 4267
rect 4456 4221 4856 4235
rect 3300 4171 3700 4185
rect 3300 4139 3334 4171
rect 3666 4139 3700 4171
rect 3300 4111 3700 4139
rect 3878 4171 4278 4185
rect 3878 4139 3902 4171
rect 4244 4139 4278 4171
rect 3878 4111 4278 4139
rect 4456 4171 4856 4185
rect 4456 4139 4678 4171
rect 4832 4139 4856 4171
rect 4456 4111 4856 4139
rect 3300 3883 3700 3911
rect 3300 3851 3334 3883
rect 3666 3851 3700 3883
rect 3300 3837 3700 3851
rect 3878 3883 4278 3911
rect 3878 3851 3902 3883
rect 4264 3851 4278 3883
rect 3878 3837 4278 3851
rect 4456 3883 4856 3911
rect 4456 3851 4678 3883
rect 4832 3851 4856 3883
rect 4456 3837 4856 3851
rect 3300 3787 3700 3801
rect 3300 3755 3324 3787
rect 3686 3755 3700 3787
rect 3300 3727 3700 3755
rect 3878 3787 4278 3801
rect 3878 3755 3902 3787
rect 4264 3755 4278 3787
rect 3878 3727 4278 3755
rect 4456 3787 4856 3801
rect 4456 3755 4470 3787
rect 4832 3755 4856 3787
rect 4456 3727 4856 3755
rect 3300 3499 3700 3527
rect 3300 3467 3324 3499
rect 3686 3467 3700 3499
rect 3300 3453 3700 3467
rect 3878 3499 4278 3527
rect 3878 3467 3892 3499
rect 4264 3467 4278 3499
rect 3878 3453 4278 3467
rect 4456 3499 4856 3527
rect 4456 3467 4470 3499
rect 4842 3467 4856 3499
rect 4456 3453 4856 3467
rect 5470 5227 5870 5273
rect 5470 4999 5870 5027
rect 5470 4967 5492 4999
rect 5852 4967 5870 4999
rect 5470 4939 5870 4967
rect 5470 4711 5870 4739
rect 5470 4679 5492 4711
rect 5852 4679 5870 4711
rect 5470 4651 5870 4679
rect 5470 4423 5870 4451
rect 5470 4391 5492 4423
rect 5852 4391 5870 4423
rect 5470 4363 5870 4391
rect 5470 4135 5870 4163
rect 5470 4103 5492 4135
rect 5852 4103 5870 4135
rect 5470 4075 5870 4103
rect 5470 3847 5870 3875
rect 5470 3815 5492 3847
rect 5852 3815 5870 3847
rect 5470 3787 5870 3815
rect 5470 3541 5870 3587
rect 3458 2992 3548 3006
rect 3458 2960 3490 2992
rect 3522 2960 3548 2992
rect 3458 2932 3548 2960
rect 3734 2992 3824 3006
rect 3734 2960 3766 2992
rect 3798 2960 3824 2992
rect 3734 2932 3824 2960
rect 3458 2842 3548 2872
rect 3458 2810 3490 2842
rect 3522 2810 3548 2842
rect 3458 2794 3548 2810
rect 3734 2840 3824 2872
rect 3734 2808 3766 2840
rect 3798 2808 3824 2840
rect 3734 2794 3824 2808
rect 3476 2354 3556 2368
rect 3476 2322 3502 2354
rect 3534 2322 3556 2354
rect 3476 2294 3556 2322
rect 3734 2354 3814 2368
rect 3734 2322 3760 2354
rect 3792 2322 3814 2354
rect 3734 2294 3814 2322
rect 3476 2206 3556 2234
rect 3476 2174 3502 2206
rect 3534 2174 3556 2206
rect 3476 2160 3556 2174
rect 3734 2206 3814 2234
rect 3734 2174 3760 2206
rect 3792 2174 3814 2206
rect 3734 2160 3814 2174
rect 3356 770 3402 850
rect 3802 826 3944 850
rect 3802 794 3830 826
rect 3862 794 3898 826
rect 3930 794 3944 826
rect 3802 770 3944 794
rect 3356 614 3402 694
rect 3802 670 3944 694
rect 3802 638 3830 670
rect 3862 638 3898 670
rect 3930 638 3944 670
rect 3802 614 3944 638
rect 3356 458 3402 538
rect 3802 514 3944 538
rect 3802 482 3830 514
rect 3862 482 3898 514
rect 3930 482 3944 514
rect 3802 458 3944 482
rect 3356 302 3402 382
rect 3802 358 3944 382
rect 3802 326 3830 358
rect 3862 326 3898 358
rect 3930 326 3944 358
rect 3802 302 3944 326
rect 4332 2352 4412 2376
rect 4332 2320 4356 2352
rect 4388 2320 4412 2352
rect 4332 2292 4412 2320
rect 4488 2352 4568 2376
rect 4488 2320 4512 2352
rect 4544 2320 4568 2352
rect 4488 2292 4568 2320
rect 4644 2352 4724 2376
rect 4644 2320 4668 2352
rect 4700 2320 4724 2352
rect 4644 2292 4724 2320
rect 4800 2352 4880 2376
rect 4800 2320 4824 2352
rect 4856 2320 4880 2352
rect 4800 2292 4880 2320
rect 4956 2352 5036 2376
rect 4956 2320 4980 2352
rect 5012 2320 5036 2352
rect 4956 2292 5036 2320
rect 5112 2352 5192 2376
rect 5112 2320 5136 2352
rect 5168 2320 5192 2352
rect 5112 2292 5192 2320
rect 5268 2352 5348 2376
rect 5268 2320 5292 2352
rect 5324 2320 5348 2352
rect 5268 2292 5348 2320
rect 5424 2352 5504 2376
rect 5424 2320 5448 2352
rect 5480 2320 5504 2352
rect 5424 2292 5504 2320
rect 5580 2352 5660 2376
rect 5580 2320 5604 2352
rect 5636 2320 5660 2352
rect 5580 2292 5660 2320
rect 5736 2352 5816 2376
rect 5736 2320 5760 2352
rect 5792 2320 5816 2352
rect 5736 2292 5816 2320
rect 4332 264 4412 292
rect 4332 232 4356 264
rect 4388 232 4412 264
rect 4332 218 4412 232
rect 4488 264 4568 292
rect 4488 232 4512 264
rect 4544 232 4568 264
rect 4488 218 4568 232
rect 4644 264 4724 292
rect 4644 232 4668 264
rect 4700 232 4724 264
rect 4644 218 4724 232
rect 4800 264 4880 292
rect 4800 232 4824 264
rect 4856 232 4880 264
rect 4800 218 4880 232
rect 4956 264 5036 292
rect 4956 232 4980 264
rect 5012 232 5036 264
rect 4956 218 5036 232
rect 5112 264 5192 292
rect 5112 232 5136 264
rect 5168 232 5192 264
rect 5112 218 5192 232
rect 5268 264 5348 292
rect 5268 232 5292 264
rect 5324 232 5348 264
rect 5268 218 5348 232
rect 5424 264 5504 292
rect 5424 232 5448 264
rect 5480 232 5504 264
rect 5424 218 5504 232
rect 5580 264 5660 292
rect 5580 232 5604 264
rect 5636 232 5660 264
rect 5580 218 5660 232
rect 5736 264 5816 292
rect 5736 232 5760 264
rect 5792 232 5816 264
rect 5736 218 5816 232
<< polycont >>
rect 140 5311 212 5343
rect 140 2799 212 2831
rect 300 5311 372 5343
rect 300 2799 372 2831
rect 460 5311 532 5343
rect 460 2799 532 2831
rect 620 5311 692 5343
rect 620 2799 692 2831
rect 780 5311 852 5343
rect 780 2799 852 2831
rect 940 5311 1012 5343
rect 940 2799 1012 2831
rect 1100 5311 1172 5343
rect 1100 2799 1172 2831
rect 1260 5311 1332 5343
rect 1260 2799 1332 2831
rect 1420 5311 1492 5343
rect 1420 2799 1492 2831
rect 1580 5311 1652 5343
rect 1580 2799 1652 2831
rect 1740 5311 1812 5343
rect 1740 2799 1812 2831
rect 1900 5311 1972 5343
rect 1900 2799 1972 2831
rect 2060 5311 2132 5343
rect 2060 2799 2132 2831
rect 2220 5311 2292 5343
rect 2220 2799 2292 2831
rect 2380 5311 2452 5343
rect 2380 2799 2452 2831
rect 2540 5311 2612 5343
rect 2540 2799 2612 2831
rect 2700 5311 2772 5343
rect 2700 2799 2772 2831
rect 2858 5311 2930 5343
rect 2858 2799 2930 2831
rect 140 2615 212 2647
rect 140 103 212 135
rect 300 2615 372 2647
rect 300 103 372 135
rect 460 2615 532 2647
rect 460 103 532 135
rect 620 2615 692 2647
rect 620 103 692 135
rect 780 2615 852 2647
rect 780 103 852 135
rect 940 2615 1012 2647
rect 940 103 1012 135
rect 1100 2615 1172 2647
rect 1100 103 1172 135
rect 1260 2615 1332 2647
rect 1260 103 1332 135
rect 1420 2615 1492 2647
rect 1420 103 1492 135
rect 1580 2615 1652 2647
rect 1580 103 1652 135
rect 1740 2615 1812 2647
rect 1740 103 1812 135
rect 1900 2615 1972 2647
rect 1900 103 1972 135
rect 2060 2615 2132 2647
rect 2060 103 2132 135
rect 2220 2615 2292 2647
rect 2220 103 2292 135
rect 2380 2615 2452 2647
rect 2380 103 2452 135
rect 2540 2615 2612 2647
rect 2540 103 2612 135
rect 2700 2615 2772 2647
rect 2700 103 2772 135
rect 2858 2615 2930 2647
rect 2858 103 2930 135
rect 3324 5291 3686 5323
rect 3902 5291 4264 5323
rect 4470 5291 4832 5323
rect 3324 5003 3686 5035
rect 3902 5003 4264 5035
rect 4470 5003 4832 5035
rect 3334 4907 3666 4939
rect 3902 4907 4056 4939
rect 4470 4907 4832 4939
rect 3334 4619 3666 4651
rect 3902 4619 4056 4651
rect 4490 4619 4832 4651
rect 3334 4523 3666 4555
rect 4100 4523 4254 4555
rect 4480 4523 4634 4555
rect 3334 4235 3666 4267
rect 4100 4235 4254 4267
rect 4480 4235 4634 4267
rect 3334 4139 3666 4171
rect 3902 4139 4244 4171
rect 4678 4139 4832 4171
rect 3334 3851 3666 3883
rect 3902 3851 4264 3883
rect 4678 3851 4832 3883
rect 3324 3755 3686 3787
rect 3902 3755 4264 3787
rect 4470 3755 4832 3787
rect 3324 3467 3686 3499
rect 3892 3467 4264 3499
rect 4470 3467 4842 3499
rect 5492 4967 5852 4999
rect 5492 4679 5852 4711
rect 5492 4391 5852 4423
rect 5492 4103 5852 4135
rect 5492 3815 5852 3847
rect 3490 2960 3522 2992
rect 3766 2960 3798 2992
rect 3490 2810 3522 2842
rect 3766 2808 3798 2840
rect 3502 2322 3534 2354
rect 3760 2322 3792 2354
rect 3502 2174 3534 2206
rect 3760 2174 3792 2206
rect 3830 794 3862 826
rect 3898 794 3930 826
rect 3830 638 3862 670
rect 3898 638 3930 670
rect 3830 482 3862 514
rect 3898 482 3930 514
rect 3830 326 3862 358
rect 3898 326 3930 358
rect 4356 2320 4388 2352
rect 4512 2320 4544 2352
rect 4668 2320 4700 2352
rect 4824 2320 4856 2352
rect 4980 2320 5012 2352
rect 5136 2320 5168 2352
rect 5292 2320 5324 2352
rect 5448 2320 5480 2352
rect 5604 2320 5636 2352
rect 5760 2320 5792 2352
rect 4356 232 4388 264
rect 4512 232 4544 264
rect 4668 232 4700 264
rect 4824 232 4856 264
rect 4980 232 5012 264
rect 5136 232 5168 264
rect 5292 232 5324 264
rect 5448 232 5480 264
rect 5604 232 5636 264
rect 5760 232 5792 264
<< xpolyres >>
rect 126 2871 226 5271
rect 286 2871 386 5271
rect 446 2871 546 5271
rect 606 2871 706 5271
rect 766 2871 866 5271
rect 926 2871 1026 5271
rect 1086 2871 1186 5271
rect 1246 2871 1346 5271
rect 1406 2871 1506 5271
rect 1566 2871 1666 5271
rect 1726 2871 1826 5271
rect 1886 2871 1986 5271
rect 2046 2871 2146 5271
rect 2206 2871 2306 5271
rect 2366 2871 2466 5271
rect 2526 2871 2626 5271
rect 2686 2871 2786 5271
rect 2844 2871 2944 5271
rect 126 175 226 2575
rect 286 175 386 2575
rect 446 175 546 2575
rect 606 175 706 2575
rect 766 175 866 2575
rect 926 175 1026 2575
rect 1086 175 1186 2575
rect 1246 175 1346 2575
rect 1406 175 1506 2575
rect 1566 175 1666 2575
rect 1726 175 1826 2575
rect 1886 175 1986 2575
rect 2046 175 2146 2575
rect 2206 175 2306 2575
rect 2366 175 2466 2575
rect 2526 175 2626 2575
rect 2686 175 2786 2575
rect 2844 175 2944 2575
<< metal1 >>
rect -10 5444 3080 5445
rect 3132 5444 5026 5445
rect -10 5435 5026 5444
rect -10 10 0 5435
rect 32 5393 3038 5403
rect 32 5343 226 5393
rect 32 5311 140 5343
rect 212 5311 226 5343
rect 32 5301 226 5311
rect 286 5343 546 5357
rect 286 5311 300 5343
rect 372 5311 460 5343
rect 532 5311 546 5343
rect 286 5301 546 5311
rect 606 5343 866 5357
rect 606 5311 620 5343
rect 692 5311 780 5343
rect 852 5311 866 5343
rect 606 5301 866 5311
rect 926 5343 1186 5357
rect 926 5311 940 5343
rect 1012 5311 1100 5343
rect 1172 5311 1186 5343
rect 926 5301 1186 5311
rect 1246 5343 1506 5357
rect 1246 5311 1260 5343
rect 1332 5311 1420 5343
rect 1492 5311 1506 5343
rect 1246 5301 1506 5311
rect 1566 5343 1826 5357
rect 1566 5311 1580 5343
rect 1652 5311 1740 5343
rect 1812 5311 1826 5343
rect 1566 5301 1826 5311
rect 1886 5343 2146 5357
rect 1886 5311 1900 5343
rect 1972 5311 2060 5343
rect 2132 5311 2146 5343
rect 1886 5301 2146 5311
rect 2206 5343 2466 5357
rect 2206 5311 2220 5343
rect 2292 5311 2380 5343
rect 2452 5311 2466 5343
rect 2206 5301 2466 5311
rect 2526 5343 2786 5357
rect 2526 5311 2540 5343
rect 2612 5311 2700 5343
rect 2772 5311 2786 5343
rect 2526 5301 2786 5311
rect 2844 5343 3038 5393
rect 2844 5311 2858 5343
rect 2930 5311 3038 5343
rect 2844 5301 3038 5311
rect 32 5166 42 5301
rect 3028 5166 3038 5301
rect 32 3000 3038 5166
rect 32 2841 42 3000
rect 3028 2841 3038 3000
rect 32 2831 386 2841
rect 32 2799 140 2831
rect 212 2799 300 2831
rect 372 2799 386 2831
rect 32 2749 386 2799
rect 446 2831 706 2841
rect 446 2799 460 2831
rect 532 2799 620 2831
rect 692 2799 706 2831
rect 446 2785 706 2799
rect 766 2831 1026 2841
rect 766 2799 780 2831
rect 852 2799 940 2831
rect 1012 2799 1026 2831
rect 766 2785 1026 2799
rect 1086 2831 1346 2841
rect 1086 2799 1100 2831
rect 1172 2799 1260 2831
rect 1332 2799 1346 2831
rect 1086 2785 1346 2799
rect 1406 2831 1666 2841
rect 1406 2799 1420 2831
rect 1492 2799 1580 2831
rect 1652 2799 1666 2831
rect 1406 2785 1666 2799
rect 1726 2832 1986 2841
rect 1726 2831 1746 2832
rect 1966 2831 1986 2832
rect 1726 2799 1740 2831
rect 1972 2799 1986 2831
rect 1726 2792 1746 2799
rect 1966 2792 1986 2799
rect 1726 2785 1986 2792
rect 2046 2831 2306 2841
rect 2046 2799 2060 2831
rect 2132 2799 2220 2831
rect 2292 2799 2306 2831
rect 2046 2785 2306 2799
rect 2366 2831 2626 2841
rect 2366 2799 2380 2831
rect 2452 2799 2540 2831
rect 2612 2799 2626 2831
rect 2366 2785 2626 2799
rect 2686 2834 2786 2841
rect 2686 2794 2700 2834
rect 2772 2794 2786 2834
rect 2686 2785 2786 2794
rect 2844 2831 3038 2841
rect 2844 2799 2858 2831
rect 2930 2799 3038 2831
rect 2844 2749 3038 2799
rect 32 2697 3038 2749
rect 32 2647 226 2697
rect 32 2615 140 2647
rect 212 2615 226 2647
rect 32 2605 226 2615
rect 286 2650 546 2661
rect 286 2610 300 2650
rect 532 2610 546 2650
rect 286 2605 546 2610
rect 606 2652 866 2661
rect 606 2612 620 2652
rect 852 2612 866 2652
rect 606 2605 866 2612
rect 926 2647 1186 2661
rect 926 2615 940 2647
rect 1012 2615 1100 2647
rect 1172 2615 1186 2647
rect 926 2605 1186 2615
rect 1246 2652 1506 2661
rect 1246 2612 1260 2652
rect 1492 2612 1506 2652
rect 1246 2605 1506 2612
rect 1566 2647 1826 2661
rect 1566 2615 1580 2647
rect 1652 2615 1740 2647
rect 1812 2615 1826 2647
rect 1566 2605 1826 2615
rect 1886 2647 2146 2661
rect 1886 2615 1900 2647
rect 1972 2615 2060 2647
rect 2132 2615 2146 2647
rect 1886 2605 2146 2615
rect 2206 2647 2466 2661
rect 2206 2615 2220 2647
rect 2292 2615 2380 2647
rect 2452 2615 2466 2647
rect 2206 2605 2466 2615
rect 2526 2652 2626 2661
rect 2526 2612 2540 2652
rect 2612 2612 2626 2652
rect 2526 2605 2626 2612
rect 2686 2647 3038 2697
rect 2686 2615 2700 2647
rect 2772 2615 2858 2647
rect 2930 2615 3038 2647
rect 32 2486 42 2605
rect 2686 2486 3038 2615
rect 32 328 3038 2486
rect 32 145 42 328
rect 32 135 226 145
rect 32 103 140 135
rect 212 103 226 135
rect 32 53 226 103
rect 286 138 386 145
rect 286 98 300 138
rect 372 98 386 138
rect 286 89 386 98
rect 446 135 706 145
rect 446 103 460 135
rect 532 103 620 135
rect 692 103 706 135
rect 446 89 706 103
rect 766 135 1026 145
rect 766 103 780 135
rect 852 103 940 135
rect 1012 103 1026 135
rect 766 89 1026 103
rect 1086 135 1346 145
rect 1086 103 1100 135
rect 1172 103 1260 135
rect 1332 103 1346 135
rect 1086 89 1346 103
rect 1406 135 1666 145
rect 1406 103 1420 135
rect 1492 103 1580 135
rect 1652 103 1666 135
rect 1406 89 1666 103
rect 1726 135 1986 145
rect 1726 103 1740 135
rect 1812 103 1900 135
rect 1972 103 1986 135
rect 1726 89 1986 103
rect 2046 135 2306 145
rect 2046 103 2060 135
rect 2132 103 2220 135
rect 2292 103 2306 135
rect 2046 89 2306 103
rect 2366 135 2626 145
rect 2366 103 2380 135
rect 2452 103 2540 135
rect 2612 103 2626 135
rect 2366 89 2626 103
rect 2686 135 3038 328
rect 2686 103 2700 135
rect 2772 103 2858 135
rect 2930 103 3038 135
rect 32 52 386 53
rect 2686 52 3038 103
rect 32 42 3038 52
rect 3070 3381 3142 5435
rect 3174 5393 4984 5403
rect 3174 5249 3278 5393
rect 3314 5291 3324 5323
rect 3686 5291 3696 5323
rect 3892 5291 3902 5323
rect 4264 5295 4274 5323
rect 4460 5295 4470 5323
rect 4264 5291 4470 5295
rect 4832 5291 4842 5323
rect 3912 5249 4824 5291
rect 3174 5077 3246 5249
rect 3278 5247 3288 5249
rect 3712 5247 3722 5249
rect 3278 5079 3722 5247
rect 3278 5077 3288 5079
rect 3712 5077 3722 5079
rect 3754 5077 3764 5249
rect 3814 5077 3824 5249
rect 3856 5247 3866 5249
rect 3912 5247 4300 5249
rect 3856 5079 4300 5247
rect 3856 5077 3866 5079
rect 3912 5077 4300 5079
rect 4332 5077 4402 5249
rect 4434 5247 4824 5249
rect 4868 5247 4878 5249
rect 4434 5079 4878 5247
rect 4434 5077 4824 5079
rect 4868 5077 4878 5079
rect 4910 5077 4920 5249
rect 3174 4865 3278 5077
rect 3314 5003 3324 5035
rect 3686 5003 3696 5035
rect 3324 4939 3676 5003
rect 3324 4907 3334 4939
rect 3666 4907 3676 4939
rect 3174 4693 3246 4865
rect 3278 4693 3288 4865
rect 3174 4481 3278 4693
rect 3324 4651 3676 4907
rect 3814 4865 3856 5077
rect 3912 5035 4824 5077
rect 3892 5003 3902 5035
rect 4264 5027 4470 5035
rect 4264 5003 4274 5027
rect 4460 5003 4470 5027
rect 4832 5003 4842 5035
rect 3902 4939 4056 4949
rect 3712 4693 3722 4865
rect 3754 4693 3824 4865
rect 3856 4693 3866 4865
rect 3324 4619 3334 4651
rect 3666 4619 3676 4651
rect 3324 4555 3676 4619
rect 3324 4523 3334 4555
rect 3666 4523 3676 4555
rect 3324 4491 3676 4523
rect 3324 4481 3764 4491
rect 3174 4309 3246 4481
rect 3278 4309 3288 4481
rect 3324 4309 3722 4481
rect 3754 4309 3764 4481
rect 3174 4097 3278 4309
rect 3324 4299 3764 4309
rect 3814 4481 3856 4693
rect 3902 4651 4056 4907
rect 3814 4309 3824 4481
rect 3856 4309 3866 4481
rect 3324 4267 3676 4299
rect 3324 4235 3334 4267
rect 3666 4235 3676 4267
rect 3324 4171 3676 4235
rect 3324 4139 3334 4171
rect 3666 4139 3676 4171
rect 3174 3925 3246 4097
rect 3278 3925 3288 4097
rect 3174 3713 3278 3925
rect 3324 3883 3676 4139
rect 3814 4097 3856 4309
rect 3902 4171 4056 4619
rect 4100 4939 4832 4949
rect 4100 4928 4470 4939
rect 4100 4630 4118 4928
rect 4216 4911 4470 4928
rect 4216 4630 4254 4911
rect 4460 4907 4470 4911
rect 4100 4555 4254 4630
rect 4300 4865 4342 4875
rect 4332 4693 4342 4865
rect 4392 4855 4402 4865
rect 4434 4855 4444 4865
rect 4392 4703 4398 4855
rect 4438 4703 4444 4855
rect 4392 4693 4402 4703
rect 4434 4693 4444 4703
rect 4300 4617 4342 4693
rect 4480 4651 4832 4907
rect 4878 4865 4910 5077
rect 4868 4693 4878 4865
rect 4910 4693 4920 4865
rect 4480 4619 4490 4651
rect 4300 4575 4434 4617
rect 4100 4267 4254 4523
rect 4298 4481 4342 4491
rect 4298 4309 4300 4481
rect 4332 4471 4342 4481
rect 4340 4319 4342 4471
rect 4332 4309 4342 4319
rect 4298 4301 4342 4309
rect 4100 4225 4254 4235
rect 4300 4227 4342 4301
rect 4392 4489 4434 4575
rect 4480 4555 4634 4565
rect 4392 4481 4436 4489
rect 4392 4475 4402 4481
rect 4392 4323 4394 4475
rect 4392 4309 4402 4323
rect 4434 4309 4436 4481
rect 4392 4299 4436 4309
rect 4480 4267 4634 4523
rect 4300 4183 4434 4227
rect 4244 4139 4254 4171
rect 3712 3925 3722 4097
rect 3754 3925 3824 4097
rect 3856 3925 3866 4097
rect 3324 3851 3334 3883
rect 3666 3851 3676 3883
rect 3324 3787 3400 3851
rect 3494 3787 3676 3851
rect 3314 3755 3324 3787
rect 3686 3755 3696 3787
rect 3814 3713 3856 3925
rect 3902 3883 4254 4139
rect 4392 4097 4434 4183
rect 4290 3925 4300 4097
rect 4332 4087 4342 4097
rect 4340 3935 4342 4087
rect 4332 3925 4342 3935
rect 4392 3925 4402 4097
rect 4392 3915 4434 3925
rect 4264 3879 4274 3883
rect 4480 3879 4634 4235
rect 4264 3851 4634 3879
rect 3902 3841 4634 3851
rect 4678 4171 4832 4619
rect 4878 4481 4910 4693
rect 4868 4309 4878 4481
rect 4910 4309 4920 4481
rect 4678 3883 4832 4139
rect 4878 4097 4910 4309
rect 4868 3925 4878 4097
rect 4910 3925 4920 4097
rect 4678 3841 4832 3851
rect 4262 3838 4632 3841
rect 3892 3755 3902 3787
rect 4264 3767 4274 3787
rect 4460 3767 4470 3787
rect 4264 3755 4470 3767
rect 4832 3755 4842 3787
rect 3912 3713 4828 3755
rect 4878 3713 4910 3925
rect 3174 3541 3246 3713
rect 3278 3711 3288 3713
rect 3712 3711 3722 3713
rect 3278 3543 3722 3711
rect 3278 3541 3288 3543
rect 3712 3541 3722 3543
rect 3754 3541 3764 3713
rect 3814 3541 3824 3713
rect 3856 3711 3866 3713
rect 3912 3711 4300 3713
rect 3856 3543 4300 3711
rect 3856 3541 3866 3543
rect 3912 3541 4300 3543
rect 4332 3541 4402 3713
rect 4434 3711 4828 3713
rect 4868 3711 4878 3713
rect 4434 3543 4878 3711
rect 4434 3541 4828 3543
rect 4868 3541 4878 3543
rect 4910 3541 4920 3713
rect 3174 3423 3278 3541
rect 3912 3499 4828 3541
rect 3314 3467 3324 3499
rect 3686 3467 3696 3499
rect 3882 3467 3892 3499
rect 4264 3483 4470 3499
rect 4264 3467 4274 3483
rect 4460 3467 4470 3483
rect 4842 3467 4852 3499
rect 4974 3423 4984 5393
rect 3174 3413 4984 3423
rect 5016 3381 5026 5435
rect 5300 5367 6048 5377
rect 5300 3435 5310 5367
rect 5342 5325 6006 5335
rect 5342 5213 5350 5325
rect 5998 5213 6006 5325
rect 5342 5041 5416 5213
rect 5448 5041 5458 5213
rect 5892 5041 5902 5213
rect 5934 5041 6006 5213
rect 5342 3783 5350 5041
rect 5492 4999 5852 5011
rect 5492 4925 5852 4967
rect 5998 4925 6006 5041
rect 5406 4753 5416 4925
rect 5448 4921 5852 4925
rect 5520 4761 5852 4921
rect 5448 4753 5852 4761
rect 5892 4753 5902 4925
rect 5934 4753 6006 4925
rect 5492 4711 5852 4753
rect 5406 4637 5456 4647
rect 5406 4633 5416 4637
rect 5448 4633 5456 4637
rect 5406 4473 5410 4633
rect 5450 4473 5456 4633
rect 5406 4465 5416 4473
rect 5448 4465 5456 4473
rect 5406 4455 5456 4465
rect 5492 4423 5852 4679
rect 5998 4637 6006 4753
rect 5892 4465 5902 4637
rect 5934 4465 6006 4637
rect 5492 4349 5852 4391
rect 5998 4349 6006 4465
rect 5406 4177 5416 4349
rect 5448 4177 5852 4349
rect 5892 4177 5902 4349
rect 5934 4177 6006 4349
rect 5492 4135 5852 4177
rect 5406 4061 5456 4071
rect 5406 4053 5416 4061
rect 5448 4053 5456 4061
rect 5406 3893 5412 4053
rect 5452 3893 5456 4053
rect 5406 3889 5416 3893
rect 5448 3889 5456 3893
rect 5406 3879 5456 3889
rect 5492 3847 5852 4103
rect 5998 4061 6006 4177
rect 5892 3889 5902 4061
rect 5934 3889 6006 4061
rect 5492 3805 5852 3815
rect 5342 3773 5456 3783
rect 5998 3773 6006 3889
rect 5342 3601 5416 3773
rect 5448 3601 5456 3773
rect 5890 3601 5900 3773
rect 5932 3601 6006 3773
rect 5342 3591 5456 3601
rect 5342 3477 5350 3591
rect 5998 3477 6006 3601
rect 5342 3467 6006 3477
rect 6038 3435 6048 5367
rect 5300 3426 6048 3435
rect 3070 3371 5026 3381
rect 5294 3425 6048 3426
rect 3070 3090 3990 3371
rect 5294 3198 6044 3425
rect 3070 2718 3302 3090
rect 3334 3048 3948 3058
rect 3334 2760 3344 3048
rect 3490 2992 3522 3002
rect 3394 2950 3446 2960
rect 3394 2910 3400 2950
rect 3440 2910 3446 2950
rect 3394 2886 3404 2910
rect 3436 2886 3446 2910
rect 3394 2860 3446 2886
rect 3490 2856 3522 2960
rect 3570 2918 3712 3048
rect 3484 2846 3528 2856
rect 3484 2806 3486 2846
rect 3526 2806 3528 2846
rect 3484 2796 3528 2806
rect 3570 2760 3712 2886
rect 3766 2992 3798 3002
rect 3766 2856 3798 2960
rect 3836 2922 3888 2940
rect 3836 2882 3842 2922
rect 3882 2882 3888 2922
rect 3836 2860 3888 2882
rect 3752 2846 3798 2856
rect 3752 2806 3754 2846
rect 3794 2840 3798 2846
rect 3794 2806 3798 2808
rect 3752 2796 3798 2806
rect 3938 2760 3948 3048
rect 3334 2750 3948 2760
rect 3980 2718 3990 3090
rect 3070 2708 3990 2718
rect 3070 10 3080 2708
rect 4174 2452 6044 3198
rect 3310 2442 5984 2452
rect 3310 2104 3320 2442
rect 3352 2400 3950 2410
rect 3352 2128 3362 2400
rect 3502 2354 3534 2364
rect 3404 2324 3456 2336
rect 3404 2284 3410 2324
rect 3450 2284 3456 2324
rect 3404 2280 3456 2284
rect 3404 2248 3422 2280
rect 3454 2248 3456 2280
rect 3404 2222 3456 2248
rect 3502 2240 3534 2322
rect 3582 2280 3712 2400
rect 3760 2354 3792 2364
rect 3752 2336 3760 2346
rect 3792 2336 3796 2346
rect 3752 2296 3754 2336
rect 3794 2296 3796 2336
rect 3752 2286 3796 2296
rect 3496 2224 3540 2240
rect 3496 2184 3498 2224
rect 3538 2184 3540 2224
rect 3496 2174 3502 2184
rect 3534 2174 3540 2184
rect 3496 2164 3540 2174
rect 3582 2128 3712 2248
rect 3760 2206 3792 2286
rect 3838 2284 3898 2306
rect 3838 2244 3844 2284
rect 3884 2244 3898 2284
rect 3838 2222 3898 2244
rect 3760 2164 3792 2174
rect 3940 2128 3950 2400
rect 3352 2118 3950 2128
rect 3260 2086 3320 2104
rect 3982 2086 4176 2442
rect 3260 1944 4176 2086
rect 4208 2400 5942 2410
rect 3260 1126 3302 1944
rect 3260 1006 4176 1126
rect 3260 146 3270 1006
rect 3302 964 3990 974
rect 3302 188 3312 964
rect 3416 910 3788 918
rect 3414 908 3790 910
rect 3414 904 3416 908
rect 3788 904 3790 908
rect 3406 872 3416 904
rect 3788 872 3798 904
rect 3414 868 3416 872
rect 3788 868 3790 872
rect 3414 866 3790 868
rect 3416 858 3788 866
rect 3820 830 3944 838
rect 3820 826 3860 830
rect 3900 826 3944 830
rect 3820 794 3830 826
rect 3930 794 3944 826
rect 3820 790 3860 794
rect 3900 790 3944 794
rect 3820 784 3944 790
rect 3414 752 3790 762
rect 3414 748 3416 752
rect 3788 748 3790 752
rect 3406 716 3416 748
rect 3788 716 3798 748
rect 3414 712 3416 716
rect 3788 712 3790 716
rect 3414 702 3790 712
rect 3820 674 3944 682
rect 3820 670 3860 674
rect 3900 670 3944 674
rect 3820 638 3830 670
rect 3930 638 3944 670
rect 3820 634 3860 638
rect 3900 634 3944 638
rect 3820 628 3944 634
rect 3416 598 3788 606
rect 3414 596 3790 598
rect 3414 592 3416 596
rect 3788 592 3790 596
rect 3406 560 3416 592
rect 3788 560 3798 592
rect 3414 556 3416 560
rect 3788 556 3790 560
rect 3414 554 3790 556
rect 3416 546 3788 554
rect 3820 518 3944 526
rect 3820 514 3860 518
rect 3900 514 3944 518
rect 3820 482 3830 514
rect 3930 482 3944 514
rect 3820 478 3860 482
rect 3900 478 3944 482
rect 3820 472 3944 478
rect 3414 440 3790 450
rect 3414 436 3416 440
rect 3788 436 3790 440
rect 3406 404 3416 436
rect 3788 404 3798 436
rect 3414 400 3416 404
rect 3788 400 3790 404
rect 3414 390 3790 400
rect 3820 362 3944 370
rect 3820 358 3860 362
rect 3900 358 3944 362
rect 3820 326 3830 358
rect 3930 326 3944 358
rect 3820 322 3860 326
rect 3900 322 3944 326
rect 3820 316 3944 322
rect 3406 284 3798 286
rect 3406 244 3416 284
rect 3788 244 3798 284
rect 3406 242 3798 244
rect 3980 188 3990 964
rect 3302 178 3990 188
rect 4022 146 4176 1006
rect 4208 186 4218 2400
rect 4278 2268 4310 2400
rect 4356 2352 4388 2362
rect 4356 2278 4388 2320
rect 4512 2352 4544 2362
rect 4273 1937 4278 1947
rect 4350 2268 4394 2278
rect 4350 2060 4352 2268
rect 4392 2060 4394 2268
rect 4350 2050 4394 2060
rect 4434 2270 4466 2284
rect 4512 2278 4544 2320
rect 4310 1937 4315 1947
rect 4273 1131 4274 1937
rect 4314 1131 4315 1937
rect 4273 1116 4278 1131
rect 4310 1116 4315 1131
rect 4278 186 4310 312
rect 4356 264 4388 2050
rect 4429 994 4434 1007
rect 4506 2268 4550 2278
rect 4506 2060 4508 2268
rect 4548 2060 4550 2268
rect 4506 2050 4550 2060
rect 4590 2270 4622 2400
rect 4668 2352 4700 2362
rect 4668 2282 4700 2320
rect 4824 2352 4856 2362
rect 4466 994 4471 1007
rect 4429 314 4430 994
rect 4470 314 4471 994
rect 4429 301 4471 314
rect 4434 300 4466 301
rect 4356 222 4388 232
rect 4512 264 4544 2050
rect 4585 1938 4590 1947
rect 4662 2270 4706 2282
rect 4662 2062 4664 2270
rect 4704 2062 4706 2270
rect 4662 2052 4706 2062
rect 4746 2270 4778 2284
rect 4824 2282 4856 2320
rect 4622 1938 4627 1947
rect 4585 1132 4586 1938
rect 4626 1132 4627 1938
rect 4585 1116 4590 1132
rect 4512 222 4544 232
rect 4622 1116 4627 1132
rect 4590 186 4622 314
rect 4668 264 4700 2052
rect 4741 994 4746 1006
rect 4818 2270 4862 2282
rect 4818 2062 4820 2270
rect 4860 2062 4862 2270
rect 4818 2052 4862 2062
rect 4902 2270 4934 2400
rect 4980 2352 5012 2362
rect 4980 2282 5012 2320
rect 5136 2352 5168 2362
rect 4778 994 4783 1006
rect 4741 314 4742 994
rect 4782 314 4783 994
rect 4741 300 4783 314
rect 4668 222 4700 232
rect 4824 264 4856 2052
rect 4897 1937 4902 1947
rect 4974 2270 5018 2282
rect 4974 2062 4976 2270
rect 5016 2062 5018 2270
rect 4974 2052 5018 2062
rect 5058 2270 5090 2284
rect 5136 2282 5168 2320
rect 4934 1937 4939 1947
rect 4897 1131 4898 1937
rect 4938 1131 4939 1937
rect 4897 1116 4902 1131
rect 4824 222 4856 232
rect 4934 1116 4939 1131
rect 4902 186 4934 314
rect 4980 264 5012 2052
rect 5053 994 5058 1006
rect 5130 2270 5174 2282
rect 5130 2062 5132 2270
rect 5172 2062 5174 2270
rect 5130 2052 5174 2062
rect 5214 2270 5246 2400
rect 5292 2352 5324 2362
rect 5292 2282 5324 2320
rect 5448 2352 5480 2362
rect 5090 994 5095 1006
rect 5053 314 5054 994
rect 5094 314 5095 994
rect 5053 300 5095 314
rect 4980 222 5012 232
rect 5136 264 5168 2052
rect 5209 1937 5214 1947
rect 5286 2270 5330 2282
rect 5286 2062 5288 2270
rect 5328 2062 5330 2270
rect 5286 2052 5330 2062
rect 5370 2270 5402 2284
rect 5448 2282 5480 2320
rect 5246 1937 5251 1947
rect 5209 1131 5210 1937
rect 5250 1131 5251 1937
rect 5209 1116 5214 1131
rect 5136 222 5168 232
rect 5246 1116 5251 1131
rect 5214 186 5246 314
rect 5292 264 5324 2052
rect 5365 994 5370 1006
rect 5442 2270 5486 2282
rect 5442 2062 5444 2270
rect 5484 2062 5486 2270
rect 5442 2052 5486 2062
rect 5526 2270 5558 2400
rect 5604 2352 5636 2362
rect 5604 2280 5636 2320
rect 5760 2352 5792 2362
rect 5402 994 5407 1006
rect 5365 314 5366 994
rect 5406 314 5407 994
rect 5365 300 5407 314
rect 5292 222 5324 232
rect 5448 264 5480 2052
rect 5521 1936 5526 1947
rect 5598 2270 5642 2280
rect 5598 2062 5600 2270
rect 5640 2062 5642 2270
rect 5598 2050 5642 2062
rect 5682 2270 5714 2284
rect 5760 2280 5792 2320
rect 5558 1936 5563 1947
rect 5521 1130 5522 1936
rect 5562 1130 5563 1936
rect 5521 1116 5526 1130
rect 5448 222 5480 232
rect 5558 1116 5563 1130
rect 5526 186 5558 314
rect 5604 264 5636 2050
rect 5677 994 5682 1006
rect 5754 2270 5798 2280
rect 5754 2062 5756 2270
rect 5796 2062 5798 2270
rect 5754 2050 5798 2062
rect 5838 2270 5870 2400
rect 5714 994 5719 1006
rect 5677 314 5678 994
rect 5718 314 5719 994
rect 5677 300 5719 314
rect 5604 222 5636 232
rect 5760 264 5792 2050
rect 5833 1934 5838 1947
rect 5870 1934 5875 1947
rect 5833 1128 5834 1934
rect 5874 1128 5875 1934
rect 5833 1116 5838 1128
rect 5760 222 5792 232
rect 5870 1116 5875 1128
rect 5838 186 5870 314
rect 5932 186 5942 2400
rect 4208 176 5942 186
rect 3260 144 4176 146
rect 5974 144 5984 2442
rect 3260 136 5984 144
rect 4166 134 5984 136
rect -10 0 3080 10
<< via1 >>
rect 1746 2831 1966 2832
rect 1746 2799 1812 2831
rect 1812 2799 1900 2831
rect 1900 2799 1966 2831
rect 1746 2792 1966 2799
rect 2700 2831 2772 2834
rect 2700 2799 2772 2831
rect 2700 2794 2772 2799
rect 300 2647 532 2650
rect 300 2615 372 2647
rect 372 2615 460 2647
rect 460 2615 532 2647
rect 300 2610 532 2615
rect 620 2647 852 2652
rect 620 2615 692 2647
rect 692 2615 780 2647
rect 780 2615 852 2647
rect 620 2612 852 2615
rect 1260 2647 1492 2652
rect 1260 2615 1332 2647
rect 1332 2615 1420 2647
rect 1420 2615 1492 2647
rect 1260 2612 1492 2615
rect 2540 2647 2612 2652
rect 2540 2615 2612 2647
rect 2540 2612 2612 2615
rect 300 135 372 138
rect 300 103 372 135
rect 300 98 372 103
rect 4118 4630 4216 4928
rect 4398 4703 4402 4855
rect 4402 4703 4434 4855
rect 4434 4703 4438 4855
rect 4300 4319 4332 4471
rect 4332 4319 4340 4471
rect 4394 4323 4402 4475
rect 4402 4323 4434 4475
rect 3400 3851 3494 3868
rect 3400 3787 3494 3851
rect 3400 3778 3494 3787
rect 4300 3935 4332 4087
rect 4332 3935 4340 4087
rect 5416 4761 5448 4921
rect 5448 4761 5520 4921
rect 5410 4473 5416 4633
rect 5416 4473 5448 4633
rect 5448 4473 5450 4633
rect 5412 3893 5416 4053
rect 5416 3893 5448 4053
rect 5448 3893 5452 4053
rect 3400 2918 3440 2950
rect 3400 2910 3404 2918
rect 3404 2910 3436 2918
rect 3436 2910 3440 2918
rect 3486 2842 3526 2846
rect 3486 2810 3490 2842
rect 3490 2810 3522 2842
rect 3522 2810 3526 2842
rect 3486 2806 3526 2810
rect 3842 2918 3882 2922
rect 3842 2886 3846 2918
rect 3846 2886 3878 2918
rect 3878 2886 3882 2918
rect 3842 2882 3882 2886
rect 3754 2840 3794 2846
rect 3754 2808 3766 2840
rect 3766 2808 3794 2840
rect 3754 2806 3794 2808
rect 3410 2284 3450 2324
rect 3754 2322 3760 2336
rect 3760 2322 3792 2336
rect 3792 2322 3794 2336
rect 3754 2296 3794 2322
rect 3498 2206 3538 2224
rect 3498 2184 3502 2206
rect 3502 2184 3534 2206
rect 3534 2184 3538 2206
rect 3844 2280 3884 2284
rect 3844 2248 3848 2280
rect 3848 2248 3880 2280
rect 3880 2248 3884 2280
rect 3844 2244 3884 2248
rect 3302 1126 4176 1944
rect 4176 1126 4200 1944
rect 3416 904 3788 908
rect 3416 872 3788 904
rect 3416 868 3788 872
rect 3860 826 3900 830
rect 3860 794 3862 826
rect 3862 794 3898 826
rect 3898 794 3900 826
rect 3860 790 3900 794
rect 3416 748 3788 752
rect 3416 716 3788 748
rect 3416 712 3788 716
rect 3860 670 3900 674
rect 3860 638 3862 670
rect 3862 638 3898 670
rect 3898 638 3900 670
rect 3860 634 3900 638
rect 3416 592 3788 596
rect 3416 560 3788 592
rect 3416 556 3788 560
rect 3860 514 3900 518
rect 3860 482 3862 514
rect 3862 482 3898 514
rect 3898 482 3900 514
rect 3860 478 3900 482
rect 3416 436 3788 440
rect 3416 404 3788 436
rect 3416 400 3788 404
rect 3860 358 3900 362
rect 3860 326 3862 358
rect 3862 326 3898 358
rect 3898 326 3900 358
rect 3860 322 3900 326
rect 3416 280 3788 284
rect 3416 248 3788 280
rect 3416 244 3788 248
rect 4352 2060 4392 2268
rect 4274 1131 4278 1937
rect 4278 1131 4310 1937
rect 4310 1131 4314 1937
rect 4508 2060 4548 2268
rect 4430 314 4434 994
rect 4434 314 4466 994
rect 4466 314 4470 994
rect 4664 2062 4704 2270
rect 4586 1132 4590 1938
rect 4590 1132 4622 1938
rect 4622 1132 4626 1938
rect 4820 2062 4860 2270
rect 4742 314 4746 994
rect 4746 314 4778 994
rect 4778 314 4782 994
rect 4976 2062 5016 2270
rect 4898 1131 4902 1937
rect 4902 1131 4934 1937
rect 4934 1131 4938 1937
rect 5132 2062 5172 2270
rect 5054 314 5058 994
rect 5058 314 5090 994
rect 5090 314 5094 994
rect 5288 2062 5328 2270
rect 5210 1131 5214 1937
rect 5214 1131 5246 1937
rect 5246 1131 5250 1937
rect 5444 2062 5484 2270
rect 5366 314 5370 994
rect 5370 314 5402 994
rect 5402 314 5406 994
rect 5600 2062 5640 2270
rect 5522 1130 5526 1936
rect 5526 1130 5558 1936
rect 5558 1130 5562 1936
rect 5756 2062 5796 2270
rect 5678 314 5682 994
rect 5682 314 5714 994
rect 5714 314 5718 994
rect 5834 1128 5838 1934
rect 5838 1128 5870 1934
rect 5870 1128 5874 1934
<< metal2 >>
rect 4104 4928 4244 4942
rect 4104 4820 4118 4928
rect 1794 4638 4118 4820
rect 1794 2842 1950 4638
rect 4104 4630 4118 4638
rect 4216 4630 4244 4928
rect 5402 4921 5530 4939
rect 5402 4865 5416 4921
rect 4104 4616 4244 4630
rect 4300 4855 5416 4865
rect 4300 4703 4398 4855
rect 4438 4761 5416 4855
rect 5520 4761 5530 4921
rect 4438 4703 5530 4761
rect 4300 4693 5530 4703
rect 4300 4471 4342 4693
rect 5406 4633 5500 4647
rect 4340 4319 4342 4471
rect 4300 4301 4342 4319
rect 4392 4475 4434 4489
rect 4392 4323 4394 4475
rect 4392 4097 4434 4323
rect 5406 4473 5410 4633
rect 5450 4473 5500 4633
rect 5406 4097 5500 4473
rect 4290 4087 5500 4097
rect 4290 3935 4300 4087
rect 4340 4053 5500 4087
rect 4340 3935 5412 4053
rect 4290 3925 5412 3935
rect 3390 3868 3504 3878
rect 3390 3778 3400 3868
rect 3494 3778 3504 3868
rect 3390 3768 3504 3778
rect 3390 2950 3450 3768
rect 3390 2910 3400 2950
rect 3440 2910 3450 2950
rect 4910 3264 5330 3925
rect 5406 3893 5412 3925
rect 5452 3893 5500 4053
rect 5406 3879 5500 3893
rect 3836 2922 3882 2932
rect 3836 2882 3842 2922
rect 3476 2846 3794 2856
rect 1736 2832 1978 2842
rect 1736 2792 1746 2832
rect 1966 2792 1978 2832
rect 1736 2782 1978 2792
rect 2690 2834 2781 2844
rect 2690 2794 2700 2834
rect 2772 2795 2781 2834
rect 3476 2806 3486 2846
rect 3526 2806 3754 2846
rect 3476 2796 3794 2806
rect 2772 2794 2782 2795
rect 2690 2662 2782 2794
rect 292 2650 544 2660
rect 292 2610 300 2650
rect 532 2610 544 2650
rect 292 2600 544 2610
rect 610 2652 862 2662
rect 610 2612 620 2652
rect 852 2612 862 2652
rect 610 2602 862 2612
rect 1250 2652 1502 2662
rect 2686 2661 2782 2662
rect 1250 2612 1260 2652
rect 1492 2612 1502 2652
rect 1250 2602 1502 2612
rect 2526 2652 2782 2661
rect 2526 2612 2540 2652
rect 2612 2612 2782 2652
rect 2526 2604 2782 2612
rect 391 439 450 2600
rect 711 603 773 2602
rect 1338 778 1402 2602
rect 2690 980 2782 2604
rect 3754 2336 3794 2796
rect 3400 2324 3458 2334
rect 3400 2284 3410 2324
rect 3450 2284 3458 2324
rect 3754 2286 3794 2296
rect 3836 2294 3882 2882
rect 4910 2566 4962 3264
rect 5266 2566 5330 3264
rect 3400 2274 3458 2284
rect 3836 2284 3890 2294
rect 3400 2097 3446 2274
rect 3836 2244 3844 2284
rect 3884 2244 3890 2284
rect 4910 2274 5330 2566
rect 3836 2242 3890 2244
rect 3498 2224 3890 2242
rect 3538 2184 3890 2224
rect 3498 2172 3890 2184
rect 4274 2270 5904 2274
rect 4274 2268 4664 2270
rect 4274 2097 4352 2268
rect 3400 2060 4352 2097
rect 4392 2060 4508 2268
rect 4548 2062 4664 2268
rect 4704 2062 4820 2270
rect 4860 2062 4976 2270
rect 5016 2062 5132 2270
rect 5172 2062 5288 2270
rect 5328 2062 5444 2270
rect 5484 2062 5600 2270
rect 5640 2062 5756 2270
rect 5796 2062 5904 2270
rect 4548 2060 5903 2062
rect 3400 2051 5903 2060
rect 3400 2050 3446 2051
rect 3296 1944 5982 1956
rect 3296 1126 3302 1944
rect 4200 1938 5982 1944
rect 4200 1937 4586 1938
rect 4200 1131 4274 1937
rect 4314 1132 4586 1937
rect 4626 1937 5982 1938
rect 4626 1132 4898 1937
rect 4314 1131 4898 1132
rect 4938 1131 5210 1937
rect 5250 1936 5982 1937
rect 5250 1131 5522 1936
rect 4200 1130 5522 1131
rect 5562 1934 5982 1936
rect 5562 1130 5834 1934
rect 4200 1128 5834 1130
rect 5874 1128 5982 1934
rect 4200 1126 5982 1128
rect 3296 1116 5982 1126
rect 4182 994 5984 1006
rect 2690 908 3800 980
rect 2690 888 3416 908
rect 3406 868 3416 888
rect 3788 868 3800 908
rect 3406 858 3800 868
rect 4182 896 4430 994
rect 4470 896 4742 994
rect 4782 896 5054 994
rect 5094 896 5366 994
rect 5406 896 5678 994
rect 5718 896 5984 994
rect 3850 830 3946 864
rect 3850 790 3860 830
rect 3900 790 3946 830
rect 1338 752 3796 778
rect 3850 756 3946 790
rect 1338 714 3416 752
rect 3788 714 3796 752
rect 3416 702 3788 712
rect 3850 674 3946 706
rect 3850 634 3860 674
rect 3900 634 3946 674
rect 711 596 3799 603
rect 3850 598 3946 634
rect 711 556 3416 596
rect 3788 556 3799 596
rect 711 541 3799 556
rect 3850 518 3946 552
rect 3850 478 3860 518
rect 3900 478 3946 518
rect 3416 440 3788 450
rect 3850 444 3946 478
rect 391 400 3416 439
rect 3788 400 3799 439
rect 391 380 3799 400
rect 3850 362 3946 396
rect 3850 322 3860 362
rect 3900 322 3946 362
rect 3406 284 3802 294
rect 3850 288 3946 322
rect 3406 244 3416 284
rect 3788 244 3802 284
rect 3406 240 3802 244
rect 4182 244 4270 896
rect 5886 244 5984 896
rect 4182 240 5984 244
rect 290 147 382 148
rect 3406 147 5984 240
rect 290 138 5984 147
rect 290 98 300 138
rect 372 98 5984 138
rect 290 94 5984 98
rect 290 88 382 94
<< via2 >>
rect 4962 2566 5266 3264
rect 4270 314 4430 896
rect 4430 314 4470 896
rect 4470 314 4742 896
rect 4742 314 4782 896
rect 4782 314 5054 896
rect 5054 314 5094 896
rect 5094 314 5366 896
rect 5366 314 5406 896
rect 5406 314 5678 896
rect 5678 314 5718 896
rect 5718 314 5886 896
rect 4270 244 5886 314
<< metal3 >>
rect 4898 3264 5330 3328
rect 4898 2566 4962 3264
rect 5266 2566 5330 3264
rect 4898 2502 5330 2566
rect 4206 896 5950 960
rect 4206 244 4270 896
rect 5886 244 5950 896
rect 4206 180 5950 244
<< via3 >>
rect 4962 2566 5266 3264
rect 4270 244 5886 896
<< metal4 >>
rect 4898 3264 5330 3328
rect 4898 2566 4962 3264
rect 5266 2566 5330 3264
rect 4898 2502 5330 2566
rect 4206 896 5950 960
rect 4206 244 4270 896
rect 5886 244 5950 896
rect 4206 180 5950 244
<< via4 >>
rect 4962 2566 5266 3264
rect 4270 244 5886 896
<< metal5 >>
rect 1722 3502 3962 3622
rect 1722 1502 1842 3502
rect 3842 3326 3962 3502
rect 4898 3326 5330 3328
rect 3842 3264 5330 3326
rect 3842 2566 4962 3264
rect 5266 2566 5330 3264
rect 3842 2504 5330 2566
rect 3842 1502 3962 2504
rect 4898 2502 5330 2504
rect 1722 1382 3962 1502
rect 4206 896 5950 960
rect 4206 244 4270 896
rect 5886 244 5950 896
rect 4206 180 5950 244
<< via5 >>
rect 4962 2566 5266 3264
rect 4270 244 5886 896
<< mimcapcontact >>
rect 1842 1502 3842 3502
<< metal6 >>
rect 1722 3502 3962 3622
rect 1722 1502 1842 3502
rect 3842 1532 3962 3502
rect 4898 3264 5330 3328
rect 4898 2566 4962 3264
rect 5266 2566 5330 3264
rect 4898 2502 5330 2566
rect 3842 1502 5950 1532
rect 1722 1382 5950 1502
rect 2102 896 5950 1382
rect 2102 244 4270 896
rect 5886 244 5950 896
rect 2102 164 5950 244
<< labels >>
flabel metal2 4212 126 4270 994 0 FreeSans 320 0 0 0 out
port 5 nsew
flabel metal2 3762 2602 3782 2672 0 FreeSans 320 0 0 0 en_n
port 10 nsew
flabel metal2 3850 288 3946 396 0 FreeSans 320 0 0 0 a0
port 9 nsew
flabel metal2 3850 444 3946 552 0 FreeSans 320 0 0 0 a1
port 8 nsew
flabel metal2 3850 598 3946 706 0 FreeSans 320 0 0 0 a2
port 7 nsew
flabel metal2 3850 756 3946 864 0 FreeSans 320 0 0 0 a3
port 6 nsew
flabel metal1 3324 4266 3674 4522 1 FreeSans 320 0 0 0 ibias_1u
port 4 n
flabel metal1 456 3392 856 4660 1 FreeSans 320 0 0 0 GND
port 2 n
flabel via1 3470 1188 3934 1774 0 FreeSans 320 0 0 0 VCC
port 1 nsew
flabel metal1 4262 3838 4632 3876 1 FreeSans 320 0 0 0 ref
port 3 n
flabel metal1 4366 4925 4390 4939 3 FreeSans 320 0 0 0 ldo_ota_0.fb
flabel metal1 4352 3851 4388 3871 3 FreeSans 320 0 0 0 ldo_ota_0.ref
flabel metal1 4364 5159 4368 5197 3 FreeSans 320 0 0 0 ldo_ota_0.tail
flabel hvpsubdiffcont 5002 5165 5006 5203 3 FreeSans 320 0 0 0 ldo_ota_0.VSS
flabel hvnsubdiffcont 5324 5133 5328 5171 3 FreeSans 320 0 0 0 ldo_ota_0.VCC
flabel metal1 3672 4299 3728 4491 0 FreeSans 320 0 0 0 ldo_ota_0.ibias_1u
flabel metal2 5102 3979 5140 4073 3 FreeSans 320 0 0 0 ldo_ota_0.vg
flabel metal1 1726 2785 1986 2841 1 FreeSans 320 0 0 0 ldo3v3_Rdiv_0.fb
flabel metal1 1246 2605 1506 2661 1 FreeSans 320 0 0 0 ldo3v3_Rdiv_0.four
flabel metal1 606 2605 866 2661 1 FreeSans 320 0 0 0 ldo3v3_Rdiv_0.two
flabel metal1 286 2605 546 2661 1 FreeSans 320 0 0 0 ldo3v3_Rdiv_0.one
flabel metal1 286 89 386 145 1 FreeSans 320 0 0 0 ldo3v3_Rdiv_0.out
flabel metal2 2690 2604 2700 2707 1 FreeSans 320 0 0 0 ldo3v3_Rdiv_0.eight
<< end >>
